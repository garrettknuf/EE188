----------------------------------------------------------------------------
--
--  SH-2 Control Unit
--
--  This is an implementation of 
--
--  Entities included are:
--    
--
--  Revision History:
--     18 April 2025    Garrett Knuf    Initial revision.
--
----------------------------------------------------------------------------

--
-- Package containing constants for the control unit.
--

library ieee;
use ieee.std_logic_1164.all;
use work.GenericConstants.all;
use work.RegArrayConstants.all;

package CUConstants is

    -- ALUOpASel - select input for ALUOpA
    constant ALUOpASel_RegA  : integer range 3 downto 0 := 0;   -- RegA of RegArray
    constant ALUOpASel_DB    : integer range 3 downto 0 := 1; 
    constant ALUOpASel_Zero  : integer range 3 downto 0 := 2; 

    -- ALUOpBSel - select input for ALUOpB
    constant ALUOpBSel_RegB         : integer range 5 downto 0 := 0;    -- RegB of RegArray
    constant ALUOpBSel_Imm_Signed   : integer range 5 downto 0 := 1;    -- immediate signed
    constant ALUOpBSel_Imm_Unsigned : integer range 5 downto 0 := 2;    -- immediate unsigned
    constant ALUOpBSel_Tbit         : integer range 5 downto 0 := 3;    -- t-bit

    -- RegInSel - select where to save input to RegIn
    constant RegInSelCmd_Rn : integer range 2 downto 0 := 0;    -- generic register
    constant RegInSelCmd_R0 : integer range 2 downto 0 := 1;    -- register R0
    constant RegInSelCmd_R15 : integer range 2 downto 0 := 2;    -- register R15

    -- RegASelCmd - select what RegA outputs
    constant RegASelCmd_Rn : integer range 2 downto 0 := 0;     -- generic register
    constant RegASelCmd_DB : integer range 2 downto 0 := 1;     -- databus
    constant RegASelCmd_R0 : integer range 2 downto 0 := 2;     -- register R0

    -- RegBSelCmd - select what RegB outputs
    constant RegBSelCmd_Rm : integer range 2 downto 0 := 0;     -- generic register
    constant RegBSelCmd_R0 : integer range 2 downto 0 := 1;     -- register R0
    constant RegBSelCmd_Rn : integer range 2 downto 0 := 2;     -- generic register
    
    -- RegA1SelCmd - select what RegA1 outputs
    constant RegA1SelCmd_Rn : integer range 2 downto 0 := 0;
    constant RegA1SelCmd_Rm : integer range 2 downto 0 := 1;
    constant RegA1SelCmd_R0 : integer range 2 downto 0 := 2;

    -- RegAxInSelCmd - select what RegA1 outputs
    constant RegAxInSelCmd_Rn : integer range 2 downto 0 := 0;
    constant RegAxInSelCmd_Rm : integer range 2 downto 0 := 1;
    constant RegAxInSelCmd_R0 : integer range 2 downto 0 := 2;

    -- DBOutSel - select output of databus
    constant DBOutSel_Result : integer range 5 downto 0 := 0;
    constant DBOutSel_SR     : integer range 5 downto 0 := 1;
    constant DBOutSel_GBR    : integer range 5 downto 0 := 2;
    constant DBOutSel_VBR    : integer range 5 downto 0 := 3;
    constant DBOutSel_PR     : integer range 5 downto 0 := 4;
    constant DBOutSel_PC     : integer range 5 downto 0 := 5;

    -- ABSel - select output of address bus
    constant ABOutSel_Prog : integer range 1 downto 0 := 0;
    constant ABOutSel_Data : integer range 1 downto 0 := 1;

    -- DataAccessMode - size of data access (read or write)
    constant DataAccessMode_BYTE : integer range 2 downto 0 := 0;
    constant DataAccessMode_WORD : integer range 2 downto 0 := 1;
    constant DataAccessMode_LONG : integer range 2 downto 0 := 2;

    constant DBInMode_Signed : integer range 1 downto 0 := 0;
    constant DBInMode_Unsigned : integer range 1 downto 0 := 1;

    constant TempRegSel_Offset8 : integer range 4 downto 0 := 0;
    constant TempRegSel_Offset12 : integer range 4 downto 0 := 1;
    constant TempRegSel_RegB : integer range 4 downto 0 := 2;

    constant REGAXDATAIN_CNT : integer := 6;
    constant RegAxDataIn_AddrIDOut  : integer range REGAXDATAIN_CNT-1 downto 0 := 0;
    constant RegAxDataIn_DataAddr   : integer range REGAXDATAIN_CNT-1 downto 0 := 1;
    constant RegAxDataIn_SR         : integer range REGAXDATAIN_CNT-1 downto 0 := 2;
    constant RegAxDataIn_GBR        : integer range REGAXDATAIN_CNT-1 downto 0 := 3;
    constant RegAxDataIn_VBR        : integer range REGAXDATAIN_CNT-1 downto 0 := 4;
    constant RegAxDataIn_PR         : integer range REGAXDATAIN_CNT-1 downto 0 := 5;

    constant unused : integer := 0;

end package;


--
--
--
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.GenericConstants.all;
use work.CUConstants.all;
use work.ALUConstants.all;
use work.TbitConstants.all;
use work.MemUnitConstants.all;
use work.DAUConstants.all;
use work.PAUConstants.all;
use work.RegArrayConstants.all;
use work.StatusRegConstants.all;
use work.OpcodeConstants.all;

entity CU is

    port (
        -- CU Input Signals
        CLK     : in    std_logic;
        RST     : in    std_logic;
        DB      : in    std_logic_vector(DATA_BUS_SIZE - 1 downto 0);
        SR      : in    std_logic_vector(REG_SIZE - 1 downto 0);
        AB      : in    std_logic_vector(DATA_BUS_SIZE - 1 downto 0);

        IR      : out   std_logic_vector(INST_SIZE - 1 downto 0) := x"DEAD";
        

        -- ALU Control Signals
        ALUOpASel   : out     integer range 2 downto 0 := 0;
        ALUOpBSel   : out     integer range 5 downto 0 := 0;
        FCmd        : out     std_logic_vector(3 downto 0);            
        CinCmd      : out     std_logic_vector(1 downto 0);            
        SCmd        : out     std_logic_vector(3 downto 0);            
        ALUCmd      : out     std_logic_vector(1 downto 0);
        TbitOp      : out     std_logic_vector(3 downto 0);

        -- StatusReg Control Signals
        UpdateSR    : out   std_logic;
        SRSel       : out   integer range SRSEL_CNT-1 downto 0;

        -- PAU Control Signals
        PAU_SrcSel      : out   integer range PAU_SRC_CNT - 1 downto 0;
        PAU_OffsetSel   : out   integer range PAU_OFFSET_CNT - 1 downto 0;
        PAU_UpdatePC    : out   std_logic;
        PAU_PRSel       : out   integer range PRSEL_CNT-1 downto 0;
        PAU_IncDecBit   : out   integer range 2 downto 0;
        PAU_PrePostSel  : out   std_logic;

        -- DAU Control Signals
        DAU_SrcSel      : out   integer range DAU_SRC_CNT - 1 downto 0;
        DAU_OffsetSel   : out   integer range DAU_OFFSET_CNT - 1 downto 0;
        DAU_IncDecSel   : out   std_logic;
        DAU_IncDecBit   : out   integer range 2 downto 0;
        DAU_PrePostSel  : out   std_logic;
        DAU_GBRSel      : out   integer range GBRSEL_CNT-1 downto 0;
        DAU_VBRSel      : out   integer range VBRSEL_CNT-1 downto 0;

        -- RegArray Control Signals
        RegInSelCmd     : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegStore        : out   std_logic;
        RegASelCmd      : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegBSelCmd      : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegAxInSelCmd   : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegAxStore      : out   std_logic;
        RegA1SelCmd     : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegA2SelCmd     : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegOpSel        : out   integer  range REGOp_SrcCnt - 1 downto 0;
        RegAxDataInSel  : out   integer  range REGAXDATAIN_CNT-1 downto 0;
    
        -- IO Control signals
        DBOutSel : out integer range 5 downto 0;
        ABOutSel : out integer range 1 downto 0;
        DBInMode : out integer range 1 downto 0;
        RD     : out   std_logic;
        WR     : out   std_logic;
        DataAccessMode : out integer range 2 downto 0;

        TempReg : out std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
        TempRegSel : out integer range 4 downto 0;

        RegB : in std_logic_vector(REG_SIZE - 1 downto 0)
    );

end CU;

architecture behavioral of CU is

    constant Normal             : integer := 0;
    constant WaitForFetch       : integer := 1;
    constant BranchSlot         : integer := 2;
    constant BranchSlotRet      : integer := 3;
    constant BranchSlotDirect   : integer := 4;
    constant BootReadSP         : integer := 5;
    constant BootWaitForFetch   : integer := 6;

    constant Sleep : integer := 7;
    constant STATE_CNT      : integer := 8;

    signal NextState : integer range STATE_CNT-1 downto 0;
    signal CurrentState : integer range STATE_CNT-1 downto 0;

    signal UpdateIR : std_logic;

    signal Tbit : std_logic;

    signal UpdateTempReg : std_logic;

    signal TempRegMuxOut : std_logic_vector(31 downto 0);

begin

    Tbit <= SR(0);

    --
    TempRegMuxOut <= (31 downto 9 => IR(7)) & IR(7 downto 0) & '0' when TempRegSel = TempRegSel_Offset8 else
                    (31 downto 13 => IR(11)) & IR(11 downto 0) & '0' when TempRegSel = TempRegSel_Offset12 else
                    RegB when TempRegSel = TempRegSel_RegB else
                    (others => 'X');

    -- Control Unit Registers
    process (CLK)
    begin

        if rising_edge(CLK) then
            if RST = '1' then
                -- Since databus is 32-bits, the IR is the high 16 bits when the
                -- program address when is at an address that is a multiple of 4.
                -- When it's not a multiple of 4 them the IR is the low 16 bits.
                IR <= DB(31 downto 16) when UpdateIR = '1' and AB(1 downto 0) = "00" else
                      DB(15 downto 0) when UpdateIR = '1' and AB(1 downto 0) = "10" else
                      IR;


                --
                TempReg <= TempRegMuxOut when UpdateTempReg = '1' else TempReg;

                -- Set state of FSM
                CurrentState <= NextState;
            else
                -- Reset to idle instruction (rising edge after reset)
                IR <= OpBoot;
                CurrentState <= Normal;
            end if;

        end if;
    end process;
    
    process (all)
    begin

    -- Instruction decoding (auto-generated)
    if std_match(IR, OpMOV_Imm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Signed;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_At_Disp_PC_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_At_Disp_PC_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOV_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_Rm_To_At_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_Rm_To_At_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_Rm_To_At_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_At_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_At_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_At_Rm_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_Rm_To_At_Dec_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 0;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_Rm_To_At_Dec_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 1;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_Rm_To_At_Dec_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_At_Rm_Inc_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rm;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_At_Rm_Inc_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 1;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rm;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_At_Rm_Inc_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rm;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_R0_To_At_Disp_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_R0_To_At_Disp_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_R0_To_At_Disp_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_At_Disp_Rm_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_At_Disp_Rm_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_At_Disp_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_Rm_To_At_R0_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_Rm_To_At_R0_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_Rm_To_At_R0_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_At_R0_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_At_R0_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_At_R0_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_R0_To_At_Disp_GBR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_R0_To_At_Disp_GBR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_R0_To_At_Disp_GBR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVB_At_Disp_GBR_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= ReginSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVW_At_Disp_GBR_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= ReginSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVL_At_Disp_GBR_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= ReginSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVA) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= ReginSelCmd_R0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_R0;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_DataAddr;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpMOVT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Tbit;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSwapB) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_SWAPB;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSwapW) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_SWAPW;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpXTRCT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_XTRCT;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpADD_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpADD_Imm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Signed;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpADDC) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_CIN;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpADDV) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Overflow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_EQ_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Signed;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_EQ_RmRn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_HS) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_GE) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GEQ;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_HI) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_HI;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_GT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GT;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_PL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_Zero;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_PL;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_PZ) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_Zero;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_PZ;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCMP_STR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_STR;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpDT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_ONE;
			CinCmd <= CinCmd_Zero;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpEXTS_B) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_EXTSB;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpEXTS_W) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_EXTSW;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpEXTU_B) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_EXTUB;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpEXTU_W) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_EXTUW;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpNEG) then
			ALUOpASel <= ALUOpASel_Zero;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpNEGC) then
			ALUOpASel <= ALUOpASel_Zero;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_CINBAR;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Borrow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSUB) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSUBC) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_CINBAR;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Borrow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSUBV) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Overflow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpAND_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_AND;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpAND_Imm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpAND_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '0';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpNOT) then
			ALUOpASel <= unused;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpOR_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_OR;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpOR_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_OR;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpOR_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_OR;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '0';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpTAS_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_ONE;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '0';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpTST_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_AND;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpTST_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpTST_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '0';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpXOR_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_XOR;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpXOR_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_XOR;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpXOR_Imm_B) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_XOR;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '0';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpROTL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_ROL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpROTR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_ROR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpROTCL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_RLC;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpROTCR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_RRC;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHAL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHAR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_ASR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLL2) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSL2;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLR2) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSR2;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLL8) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSL8;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLR8) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSR8;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLL16) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSL16;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpSHLR16) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= SCmd_LSR16;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBF) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when Tbit = '0' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBFS) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot when SR(0)='0' else Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset8;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBT) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when Tbit = '1' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBTS) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot when SR(0)='1' else Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset8;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBRA) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset12;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBRAF) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBSR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_PC;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset12;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpBSRF) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_PC;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpJMP) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlotDirect;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpJSR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_PC;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlotDirect;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpRTS) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlotRet;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
		elsif std_match(IR, OpCLRT) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= FCmd_ONE;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpLDC_Rm_To_SR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= SRSel_Reg;
		elsif std_match(IR, OpLDC_Rm_To_GBR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_Reg;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpLDC_Rm_To_VBR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_Reg;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_SR) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= unused;
			FCmd <= FCmd_A;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= (others => '-');
			UpdateSR <= '1';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= SRSel_DB;
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_GBR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_DB;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_VBR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_DB;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpLDS_Rm_To_PR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_Reg;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpLDSL_At_Rm_Inc_To_PR) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_DB;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSLEEP) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= 0;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Sleep;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpNOP) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpRTE) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_OffsetReg;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '0';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSETT) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= FCmd_ZERO;
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTC_SR_To_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_SR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTC_GBR_To_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_GBR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTC_VBR_To_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_VBR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTCL_SR_To_At_Dec_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_SR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTCL_GBR_To_At_Dec_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_GBR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTCL_VBR_To_At_Dec_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_VBR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTS_PR_To_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_PR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpSTSL_PR_To_At_Dec_Rn) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_PR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpTRAPA) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= unused;
			PAU_OffsetSel <= unused;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= RegOp_None;
			RegAxDataInSel <= RegAxDataIn_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		elsif std_match(IR, OpBoot) then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrDB;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_IncDecBit <= unused;
			PAU_PrePostSel <= MemUnit_POST;
			DAU_SrcSel <= DAU_AddrZero;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= 0;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegA2SelCmd <= 0;
			RegOpSel <= 0;
			RegAxDataInSel <= 0;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= BootReadSP;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
		end if;

		-- State Decoding Autogen
		if CurrentState = WaitForFetch then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= 0;
			DAU_VBRSel <= 0;
			RegInSelCmd <= unused;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = Sleep then
			ALUOpASel <= unused;
			ALUOpBSel <= unused;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= 0;
			DAU_VBRSel <= 0;
			RegInSelCmd <= unused;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RD <= '1';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Sleep;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = BranchSlot then
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_TempReg;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			NextState <= Normal;
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			PAU_IncDecBit <= 1;
			PAU_PrePostSel <= MemUnit_PRE;
		elsif CurrentState = BranchSlotRet then
			PAU_SrcSel <= PAU_AddrPR;
			PAU_OffsetSel <= PAU_OffsetLong;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			NextState <= Normal;
			UpdateTempReg <= '1';
			TempRegSel <= unused;
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = BranchSlotDirect then
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_TempReg;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			NextState <= Normal;
			UpdateTempReg <= '1';
			TempRegSel <= unused;
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = BootReadSP then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			DAU_SrcSel <= DAU_AddrZero;
			DAU_OffsetSel <= DAU_OffsetLong;
			DAU_PrePostSel <= MemUnit_POST;
			RegInSelCmd <= RegInSelCmd_R15;
			RegStore <= '1';
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= BootWaitForFetch;
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_PRE;
		elsif CurrentState = BootWaitForFetch then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= (others => '-');
			CinCmd <= (others => '-');
			SCmd <= (others => '-');
			ALUCmd <= (others => '-');
			TbitOp <= (others => '-');
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			DAU_SrcSel <= unused;
			DAU_OffsetSel <= unused;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= unused;
			DAU_PrePostSel <= '-';
			DAU_GBRSel <= 0;
			DAU_VBRSel <= 0;
			RegInSelCmd <= unused;
			RegStore <= '0';
			RegASelCmd <= unused;
			RegBSelCmd <= unused;
			RegAxInSelCmd <= unused;
			RegAxStore <= '0';
			RegA1SelCmd <= unused;
			RegA2SelCmd <= unused;
			RegOpSel <= RegOp_None;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= unused;
			DBOutSel <= unused;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= unused;
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		end if;


    -- end of auto-generated code (continue process)
        
    end process;


end behavioral;
