----------------------------------------------------------------------------
--
--  Hitachi SH-2 RISC Processor
--
--  This file contains the complete top-level structural implementation of the
--  Hitachi SH-2 RISC Processor. It includes instantations of all major components:
--  ALU, RegArray, CU, PAU, DAU, and DTU. THE SH2_CPU entity defines the interface
--  of the processor and connects its internal subsystems in a structural
--  architecture. It is used for integration and testing of the full processor
--  design. The main resource for design is the SuperH RISC Engine SH-1/SH-2
--  Progamming Manual by Hitachi September 3, 1996.
--
--  The processor contains a 5-stage pipeline. The pipeline integrates hazard
--  detection and forwarding logic for efficient instruction throughput. The 
--  stages of the pipeline are:
--   1. IF (Instruction Fetch) - Fetches an instruction from the memory in which
--      the program is stored.
--   2. ID (Instruction Decode) - Decodes the instruction fetched.
--   3. EX (Execute) - Performs data operations and address calculations according
--      to the results of the decoding
--   4. MA (Memory Access) - Access data in memory. Generated by instructions that
--      involve memory access, with some exceptions.
--   5. WB (Writeback) - Returns the results of the memory access (data) to a register.
--      Generated by instructions that involve memory loads, with some exceptions.
--
--  Entities included are:
--    SH2_CPU - top level structural of CPU
--
--  Revision History:
--     16 Apr 2025      Garrett Knuf    Initial revision.
--     22 Apr 2025      Garrett Knuf    Integrated all components together.
--     13 May 2025      Garrett Knuf    Connect DTU.
--     16 May 2025      George Ore      Make interface synthesizable.
--     2  Jun 2025      Garrett Knuf    Add pipeline stages.
--
----------------------------------------------------------------------------

--
--  SH2_CPU
--
--  This is the complete entity declaration for the SH-2 CPU.  It is used to
--  test the complete design.
--
--  Inputs:
--    Reset  - active low reset signal
--    NMI    - active falling edge non-maskable interrupt
--    INT    - active low maskable interrupt
--    clock  - the system clock
--
--  Outputs:
--    AB     - memory address bus (32 bits)
--    RE0    - first byte read signal, active low
--    RE1    - second byte read signal, active low
--    RE2    - third byte read signal, active low
--    RE3    - fourth byte read signal, active low
--    WE0    - first byte write signal, active low
--    WE1    - second byte write signal, active low
--    WE2    - third byte write signal, active low
--    WE3    - fourth byte write signal, active low
--
--  Inputs/Outputs:
--    DB     - memory data bus (32 bits)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.GenericConstants.all;
use work.GenericALUConstants.all;
use work.ALUConstants.all;
use work.GenericALUConstants.all;
use work.MemUnitConstants.all;
use work.PAUConstants.all;
use work.DAUConstants.all;
use work.RegArrayConstants.all;
use work.CUConstants.all;
use work.DTUConstants.all;

entity  SH2_CPU  is

    port (
        Reset   :  in     std_logic;                       -- reset signal (active low)
        NMI     :  in     std_logic;                       -- non-maskable interrupt signal (falling edge)
        INT     :  in     std_logic;                       -- maskable interrupt signal (active low)
        clock   :  in     std_logic;                       -- system clock
        AB      :  out    std_logic_vector(31 downto 0);   -- memory address bus
        RE0     :  out    std_logic;                       -- first byte active low read enable
        RE1     :  out    std_logic;                       -- second byte active low read enable
        RE2     :  out    std_logic;                       -- third byte active low read enable
        RE3     :  out    std_logic;                       -- fourth byte active low read enable
        WE0     :  out    std_logic;                       -- first byte active low write enable
        WE1     :  out    std_logic;                       -- second byte active low write enable
        WE2     :  out    std_logic;                       -- third byte active low write enable
        WE3     :  out    std_logic;                       -- fourth byte active low write enable
        DB      :  inout  std_logic_vector(31 downto 0)    -- memory data bus
    );

end  SH2_CPU;

architecture structural of SH2_CPU is

    component ALU is
    port (
            -- Operand inputs
            RegA     : in       std_logic_vector(LONG_SIZE - 1 downto 0);   -- RegArray RegA
            RegB     : in       std_logic_vector(LONG_SIZE - 1 downto 0);   -- RegArray RegB
            TempReg  : in       std_logic_vector(LONG_SIZE - 1 downto 0);   -- CU TempReg
            Imm      : in       std_logic_vector(IMM_SIZE - 1 downto 0);    -- Immediate value
            DBIn     : in       std_logic_vector(LONG_SIZE - 1 downto 0);   -- DataBusIn
            SR0      : in       std_logic;                                  -- StatusReg Bit0

            -- Control signals
            ALUOpASel   : in    integer range ALUOPASEL_CNT-1 downto 0;     -- operand A select
            ALUOpBSel   : in    integer range ALUOPBSEL_CNT-1 downto 0;     -- operand B select
            FCmd        : in    std_logic_vector(3 downto 0);               -- F-Block operation
            CinCmd      : in    std_logic_vector(1 downto 0);               -- carry in operation
            SCmd        : in    std_logic_vector(2 downto 0);               -- shift operation
            ALUCmd      : in    std_logic_vector(1 downto 0);               -- ALU result select
            TbitOp      : in    std_logic_vector(3 downto 0);               -- T-bit operation

            -- Outputs
            Result   : out      std_logic_vector(LONG_SIZE - 1 downto 0);   -- ALU Result
            TBit     : out      std_logic                                   -- Calculated T bit
        );
    end component;

    component RegArray is
        port (
            -- RegIn input
            Result      : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- ALU Result

            -- RegAxIn inputs
            DataAddrID  : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- DAU inc/dec address
            DataAddr    : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- DAU address
            SR          : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- Status register
            GBR         : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- Global base register
            VBR         : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- Vector base register
            PR          : in   std_logic_vector(LONG_SIZE - 1 downto 0);    -- Procedure register

            -- Control signals
            RegInSel        : in   integer range REGARRAY_RegCnt - 1 downto 0;      -- select where to save Result
            RegStore        : in   std_logic;                                       -- decide store result or not
            RegASel         : in   integer range REGARRAY_RegCnt - 1 downto 0;      -- select RegA output
            RegBSel         : in   integer range REGARRAY_RegCnt - 1 downto 0;      -- select RegB output
            RegAxInSel      : in   integer range REGARRAY_RegCnt - 1 downto 0;      -- select where to save RegAxIn input
            RegAxInDataSel  : in   integer range REGAXINDATASEL_CNT - 1 downto 0;   -- select input to RegAxIn
            RegAxStore      : in   std_logic;                                       -- decide store RegAxIn or not
            RegA1Sel        : in   integer range REGARRAY_RegCnt - 1 downto 0;      -- select RegA1 output
            RegOpSel        : in   integer range REGOPSEL_CNT - 1 downto 0;         -- select special register operation
            CLK             : in   std_logic;                                       -- system clock

            -- Register Outputs
            RegA            : out  std_logic_vector(REG_SIZE - 1 downto 0);     -- register A
            RegB            : out  std_logic_vector(REG_SIZE - 1 downto 0);     -- register B
            RegA1           : out  std_logic_vector(REG_SIZE - 1 downto 0)      -- register Addr1
        );
    end component;

    component PAU is
        port (
            -- Control signals
            SrcSel      : in    integer range PAU_SRC_CNT - 1 downto 0;         -- source select
            OffsetSel   : in    integer range PAU_OFFSET_CNT - 1 downto 0;      -- offset select
            UpdatePC    : in    std_logic;                                      -- update PC or hold
            PRSel       : in    integer range PRSEL_CNT-1 downto 0;             -- select modify PR
            IncDecSel   : in    std_logic;                                      -- select inc/dec
            IncDecBit   : in    integer range 2 downto 0;                       -- select bit to inc/dec
            PrePostSel  : in    std_logic;                                      -- select decrement by 4

            -- Source inputs
            DB          : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- data bus
            PC_EX       : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- pipelined PC (delayed by two clocks)

            -- Offset inputs
            Offset8     : in    std_logic_vector(7 downto 0);                   -- 8-bit offset
            Offset12    : in    std_logic_vector(11 downto 0);                  -- 12-bit offset
            OffsetReg   : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- register offest
            TempReg     : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- temporary register offset

            -- System signal
            CLK         : in    std_logic;                                      -- clock
            RESET       : in    std_logic;                                      -- reset

            -- Output signals
            ProgAddr    : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- program address
            PC          : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- program counter
            PR          : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0)    -- procedure register
        );
    end component;

    component DAU is
        port (
            -- Source inputs
            PC          : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- program counter
            Rn          : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- generic register

            -- Offset inputs
            Offset4     : in    std_logic_vector(3 downto 0);                   -- 4-bit offset
            Offset8     : in    std_logic_vector(7 downto 0);                   -- 8-bit offset
            R0          : in    std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- register R0

            -- Data bus input
            DB          : in    std_logic_vector(DATA_BUS_SIZE - 1 downto 0);   -- databus

            -- Control signals
            SrcSel      : in    integer range DAU_SRC_CNT - 1 downto 0;         -- source select
            OffsetSel   : in    integer range DAU_OFFSET_CNT - 1 downto 0;      -- offset select
            IncDecSel   : in    std_logic;                                      -- select inc/dec
            IncDecBit   : in    integer range 2 downto 0;                       -- select bit to inc/dec
            PrePostSel  : in    std_logic;                                      -- select pre/post
            GBRSel      : in    integer range GBRSel_CNT-1 downto 0;            -- select GBR
            VBRSel      : in    integer range VBRSel_CNT-1 downto 0;            -- select VBR
            CLK         : in    std_logic;                                      -- system clock
            RST         : in    std_logic;                                      -- system reset

            -- Output signals
            AddrIDOut   : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- inc/dec address output
            DataAddr    : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- data address
            GBR         : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);   -- global base register
            VBR         : out   std_logic_vector(ADDR_BUS_SIZE - 1 downto 0)    -- vector base register
        );
    end component;

    component CU is
        port (
            -- CU Input Signals
            CLK     : in    std_logic;                                      -- system clock
            RST     : in    std_logic;                                      -- system reset
            DB      : in    std_logic_vector(DATA_BUS_SIZE - 1 downto 0);   -- data bus
            AB      : in    std_logic_vector(1 downto 0);                   -- address bus (least 2 significant bits)
            Result  : in    std_logic_vector(LONG_SIZE - 1 downto 0);       -- ALU result
            Tbit    : in    std_logic;                                      -- Tbit from ALU
            RegB    : in    std_logic_vector(REG_SIZE - 1 downto 0);

            -- CU Registers
            IR      : out   std_logic_vector(INST_SIZE - 1 downto 0) := x"DEAD";    -- instruction register
            SR      : out std_logic_vector(REG_SIZE - 1 downto 0);                  -- status register
            TempReg : out std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);             -- temporary register
            TempReg2 : out std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);            -- secondary temp register
            
            -- CU Output Signals
            UpdateIR    : out   std_logic;  -- update instruction register (ID stage)
            UpdateIR_EX : in std_logic;     -- pipelined signal to update IR (used to detect memory access)
            UpdateSR    : out   std_logic;  -- update status register (ID stage)
            UpdateSR_EX : in std_logic;     -- pipelined signal to update SR (used to determine conditional branching)
            SRSel       : out integer range SRSEL_CNT-1 downto 0; -- select input to status register
            SRSel_EX    : in  integer range SRSEL_CNT-1 downto 0; -- select input to status register
            
            -- ALU Control Signals
            ALUOpASel   : out     integer range ALUOPASEL_CNT-1 downto 0 := 0;  -- select operand A
            ALUOpBSel   : out     integer range ALUOPBSEL_CNT-1 downto 0 := 0;  -- select operand B
            FCmd        : out     std_logic_vector(3 downto 0);                 -- Fblock control
            CinCmd      : out     std_logic_vector(1 downto 0);                 -- carry in
            SCmd        : out     std_logic_vector(2 downto 0);                 -- shift block control
            ALUCmd      : out     std_logic_vector(1 downto 0);                 -- output mux
            TbitOp      : out     std_logic_vector(3 downto 0);                 -- tbit control

            -- PAU Control Signals
            PAU_SrcSel      : out   integer range PAU_SRC_CNT - 1 downto 0;     -- select address source
            PAU_OffsetSel   : out   integer range PAU_OFFSET_CNT - 1 downto 0;  -- select offset source
            PAU_UpdatePC    : out   std_logic;                                  -- update PC
            PAU_PRSel       : out   integer range PRSEL_CNT-1 downto 0;         -- select PR control
            PAU_IncDecSel   : out   std_logic;                                  -- select for inc/dec
            PAU_IncDecBit   : out   integer range 2 downto 0;                   -- select inc/dec
            PAU_PrePostSel  : out   std_logic;                                  -- select pre/post

            -- DAU Control Signals
            DAU_SrcSel      : out   integer range DAU_SRC_CNT - 1 downto 0;     -- select address source
            DAU_OffsetSel   : out   integer range DAU_OFFSET_CNT - 1 downto 0;  -- select offset source
            DAU_IncDecSel   : out   std_logic;                                  -- select inc/dec
            DAU_IncDecBit   : out   integer range 2 downto 0;                   -- select inc/dec bit
            DAU_PrePostSel  : out   std_logic;                                  -- select pre/post
            DAU_GBRSel      : out   integer range GBRSEL_CNT-1 downto 0;        -- select GBR load
            DAU_VBRSel      : out   integer range VBRSEL_CNT-1 downto 0;        -- select VBR load

            -- RegArray Control Signals
            RegInSel        : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select input reg
            RegStore        : out   std_logic;                                      -- store input reg
            RegASel         : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select output RegA
            RegBSel         : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select output regB
            RegAxInSel      : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select address input reg
            RegAxInDataSel  : out   integer range REGAXINDATASEL_CNT - 1 downto 0;  -- select data to address input
            RegAxStore      : out   std_logic;                                      -- store address input
            RegA1Sel        : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select address reg output
            RegOpSel        : out   integer  range REGOPSEL_CNT - 1 downto 0;       -- select special reg operation
        
            -- IO Control signals
            DBOutSel : out integer range DBOUTSEL_CNT-1 downto 0;   -- select databus output
            ABOutSel : out integer range 1 downto 0;                -- select addressbus output
            DBInMode : out integer range 1 downto 0;                -- select sign/unsigned databus read
            RD     : out   std_logic;                               -- read (active-low)
            WR     : out   std_logic;                               -- write (active-low)
            DataAccessMode : out integer range 2 downto 0;          -- align bytes, words, long

            -- Pipeline control signals
            StallPL         : out std_logic;    -- used to indicate when a pipeline stall is needed
            TakeBranch      : in std_logic;    -- used to override the next state to normal when flushing pipeline
            RMW             : out std_logic;    -- high when there is a read-modify-write (RMW) instruction
            UseWB           : out std_logic;   -- used to determine when the write back state is used
            BranchSel       : out integer range BRANCHSEL_CNT-1 downto 0  -- used to select type of branch (if any)
        );
    end component;

    component DTU is
        port (
            -- Data input
            DBOut           : in    std_logic_vector(DATA_BUS_SIZE-1 downto 0);     -- data to output to DB

            -- Control inputs
            AB              : in    std_logic_vector(1 downto 0);                   -- address bus (least 2 significant bits)
            RD              : in    std_logic;                                      -- read enable (active-low)
            WR              : in    std_logic;                                      -- write enable (active-low)
            DataAccessMode  : in    integer range DATAACCESSMODE_CNT-1 downto 0;    -- select byte, word, long access
            DBInMode        : in    integer range DBINMODE_CNT-1 downto 0;          -- select signed or unsigned read
            CLK             : in    std_logic;                                      -- system clock

            -- Control outputs
            DBIn            : out   std_logic_vector(DATA_BUS_SIZE-1 downto 0);     -- data read from DB
            WE0             : out   std_logic;                                      -- write enable byte0
            WE1             : out   std_logic;                                      -- write enable byte1
            WE2             : out   std_logic;                                      -- write enable byte2
            WE3             : out   std_logic;                                      -- write enable byte3
            RE0             : out   std_logic;                                      -- read enable byte0
            RE1             : out   std_logic;                                      -- read enable byte1
            RE2             : out   std_logic;                                      -- read enable byte2
            RE3             : out   std_logic;                                      -- read enable byte3

            -- In/Out data bus
            DB              : inout std_logic_vector(DATA_BUS_SIZE-1 downto 0)      -- data bus
        );
    end component;

    ---------------------------------------------------------------------------
    -- ALU Signals
    ---------------------------------------------------------------------------

    -- ALU ID Stage (CU -> DFFs)
    signal ALUOpASel_ID    : integer range ALUOPASEL_CNT-1 downto 0;
    signal ALUOpBSel_ID    : integer range ALUOPBSEL_CNT-1 downto 0;
    signal ALU_FCmd_ID     : std_logic_vector(3 downto 0);
    signal ALU_CinCmd_ID   : std_logic_vector(1 downto 0);
    signal ALU_SCmd_ID     : std_logic_vector(2 downto 0);
    signal ALU_ALUCmd_ID   : std_logic_vector(1 downto 0);
    signal ALU_TbitOp_ID   : std_logic_vector(3 downto 0);

    -- ALU EX Stage (DFFs -> ALU)
    signal ALUOpASel_EX    : integer range ALUOPASEL_CNT-1 downto 0;
    signal ALUOpBSel_EX    : integer range ALUOPBSEL_CNT-1 downto 0;
    signal ALU_FCmd_EX     : std_logic_vector(3 downto 0);
    signal ALU_CinCmd_EX   : std_logic_vector(1 downto 0);
    signal ALU_SCmd_EX     : std_logic_vector(2 downto 0);
    signal ALU_ALUCmd_EX   : std_logic_vector(1 downto 0);
    signal ALU_TbitOp_EX   : std_logic_vector(3 downto 0);

    -- Non-pipelined outputs
    signal ALU_Result    : std_logic_vector(LONG_SIZE - 1 downto 0);
    signal ALU_Tbit      : std_logic;

    ---------------------------------------------------------------------------
    -- RegArray Signals
    ---------------------------------------------------------------------------

    -- RegArray ID Stage (CU -> DFFs)
    signal RegInSel_ID   : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegStore_ID   : std_logic;
    signal RegASel_ID    : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegBSel_ID    : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInSel_ID : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInDataSel_ID : integer range REGAXINDATASEL_CNT - 1 downto 0;
    signal RegAxStore_ID : std_logic;
    signal RegA1Sel_ID   : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegOpSel_ID   : integer range REGOPSEL_CNT - 1 downto 0;

    -- RegArray EX Stage (DFFs -> DFFs/RegArray)
    signal RegInSel_EX   : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegStore_EX   : std_logic;
    signal RegASel_EX    : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegBSel_EX    : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInSel_EX : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInDataSel_EX : integer range REGAXINDATASEL_CNT - 1 downto 0;
    signal RegAxStore_EX : std_logic;
    signal RegA1Sel_EX   : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegOpSel_EX   : integer range REGOPSEL_CNT - 1 downto 0;

    -- RegArray MA Stage (DFFs -> DFFs/RegArray)
    signal RegInSel_MA   : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegStore_MA   : std_logic;
    signal RegASel_MA    : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegBSel_MA    : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInSel_MA : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInDataSel_MA : integer range REGAXINDATASEL_CNT - 1 downto 0;
    signal RegAxStore_MA : std_logic;
    signal RegA1Sel_MA   : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegOpSel_MA   : integer range REGOPSEL_CNT - 1 downto 0;

    -- RegArray WB Stage (DFFs -> RegArray)
    signal RegInSel_WB          : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegStore_WB          : std_logic;
    signal RegAxInSel_WB        : integer range REGARRAY_RegCnt - 1 downto 0;
    signal RegAxInDataSel_WB    : integer range REGAXINDATASEL_CNT - 1 downto 0;
    signal RegAxStore_WB        : std_logic;

    -- Non-pipelined outputs
    signal RegA       : std_logic_vector(LONG_SIZE - 1 downto 0);
    signal RegB       : std_logic_vector(LONG_SIZE - 1 downto 0);
    signal RegA1      : std_logic_vector(LONG_SIZE - 1 downto 0);
    signal RegIn      : std_logic_vector(LONG_SIZE - 1 downto 0);
    signal RegAxIn    : std_logic_vector(LONG_SIZE - 1 downto 0);

    ---------------------------------------------------------------------------
    -- PAU Signals
    ---------------------------------------------------------------------------

    -- PAU ID Stage (CU -> DFFs)
    signal PAU_SrcSel_ID      : integer range PAU_SRC_CNT - 1 downto 0;
    signal PAU_OffsetSel_ID   : integer range PAU_OFFSET_CNT - 1 downto 0;
    signal PAU_UpdatePC_ID    : std_logic;
    signal PAU_PRSel_ID       : integer range PRSEL_CNT-1 downto 0;
    signal PAU_IncDecSel_ID   : std_logic;
    signal PAU_IncDecBit_ID   : integer range 2 downto 0;
    signal PAU_PrePostSel_ID  : std_logic;
    signal PC_ID              : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);

    -- PAU EX Stage (DFFs -> PAU)
    signal PAU_SrcSel_EX      : integer range PAU_SRC_CNT - 1 downto 0;
    signal PAU_OffsetSel_EX   : integer range PAU_OFFSET_CNT - 1 downto 0;
    signal PAU_UpdatePC_EX    : std_logic;
    signal PAU_PRSel_EX       : integer range PRSEL_CNT-1 downto 0;
    signal PAU_IncDecSel_EX   : std_logic;
    signal PAU_IncDecBit_EX   : integer range 2 downto 0;
    signal PAU_PrePostSel_EX  : std_logic;
    signal PC_EX              : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);

    -- Non-pipelined outputs
    signal PAU_ProgAddr    : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal PAU_OffsetReg   : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal PR              : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);

    ---------------------------------------------------------------------------
    -- DAU Signals
    ---------------------------------------------------------------------------

    -- DAU ID Stage (CU -> DFFs)
    signal DAU_SrcSel_ID      : integer range DAU_SRC_CNT - 1 downto 0;
    signal DAU_OffsetSel_ID   : integer range DAU_OFFSET_CNT - 1 downto 0;
    signal DAU_Offset4_ID     : std_logic_vector(3 downto 0);
    signal DAU_Offset8_ID     : std_logic_vector(7 downto 0);
    signal DAU_IncDecSel_ID   : std_logic;
    signal DAU_IncDecBit_ID   : integer range 2 downto 0;
    signal DAU_PrePostSel_ID  : std_logic;
    signal DAU_GBRSel_ID      : integer range GBRSEL_CNT-1 downto 0;
    signal DAU_VBRSel_ID      : integer range VBRSEL_CNT-1 downto 0;

    -- DAU EX Stage (DFFs -> DFFs/DAU)
    signal DAU_SrcSel_EX      : integer range DAU_SRC_CNT - 1 downto 0;
    signal DAU_OffsetSel_EX   : integer range DAU_OFFSET_CNT - 1 downto 0;
    signal DAU_Offset4_EX     : std_logic_vector(3 downto 0);
    signal DAU_Offset8_EX     : std_logic_vector(7 downto 0);
    signal DAU_IncDecSel_EX   : std_logic;
    signal DAU_IncDecBit_EX   : integer range 2 downto 0;
    signal DAU_PrePostSel_EX  : std_logic;
    signal DAU_GBRSel_EX      : integer range GBRSEL_CNT-1 downto 0;
    signal DAU_VBRSel_EX      : integer range VBRSEL_CNT-1 downto 0;

    -- DAU MA Stage (DFFs -> DFFs/DAU)
    signal DAU_SrcSel_MA      : integer range DAU_SRC_CNT - 1 downto 0;
    signal DAU_OffsetSel_MA   : integer range DAU_OFFSET_CNT - 1 downto 0;
    signal DAU_Offset4_MA     : std_logic_vector(3 downto 0);
    signal DAU_Offset8_MA     : std_logic_vector(7 downto 0);
    signal DAU_IncDecSel_MA   : std_logic;
    signal DAU_IncDecBit_MA   : integer range 2 downto 0;
    signal DAU_PrePostSel_MA  : std_logic;
    signal DAU_GBRSel_MA      : integer range GBRSEL_CNT-1 downto 0;
    signal DAU_VBRSel_MA      : integer range VBRSEL_CNT-1 downto 0;

    -- DAU WB Stage (DFFs -> DAU)
    signal DAU_SrcSel_WB      : integer range DAU_SRC_CNT - 1 downto 0;
    signal DAU_OffsetSel_WB   : integer range DAU_OFFSET_CNT - 1 downto 0;
    signal DAU_Offset4_WB     : std_logic_vector(3 downto 0);
    signal DAU_Offset8_WB     : std_logic_vector(7 downto 0);
    signal DAU_IncDecSel_WB   : std_logic;
    signal DAU_IncDecBit_WB   : integer range 2 downto 0;
    signal DAU_PrePostSel_WB  : std_logic;
    signal DAU_GBRSel_WB      : integer range GBRSEL_CNT-1 downto 0;
    signal DAU_VBRSel_WB      : integer range VBRSEL_CNT-1 downto 0;
    
    -- Non-pipelined outputs
    signal DAU_Rn          : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal DAU_R0          : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal DAU_PC          : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal DAU_IncDecSel   : std_logic;
    signal DAU_IncDecBit   : integer range 2 downto 0;
    signal DAU_PrePostSel  : std_logic;
    signal DAU_GBRSel      : integer range GBRSEL_CNT-1 downto 0;
    signal DAU_VBRSel      : integer range VBRSEL_CNT-1 downto 0;
    signal DAU_AddrIDOut   : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal DAU_DataAddr    : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal GBR             : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);
    signal VBR             : std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);

    ---------------------------------------------------------------------------
    -- DTU Signals
    ---------------------------------------------------------------------------

    -- DTU ID Stage (CU -> DFFs)
    signal DBInMode_ID          : integer range DBINMODE_CNT-1 downto 0;
    signal DataAccessMode_ID    : integer range DATAACCESSMODE_CNT-1 downto 0;
    signal WR_ID                : std_logic;
    signal RD_ID                : std_logic;
    
    -- DTU EX Stage (DFFs -> DFFs)
    signal DBInMode_EX          : integer range DBINMODE_CNT-1 downto 0;
    signal DataAccessMode_EX    : integer range DATAACCESSMODE_CNT-1 downto 0;
    signal WR_EX                : std_logic;
    signal RD_EX                : std_logic;

    -- DTU MA Stage (DFFs -> DFFs)
    signal DBInMode_MA          : integer range DBINMODE_CNT-1 downto 0;
    signal DataAccessMode_MA    : integer range DATAACCESSMODE_CNT-1 downto 0;
    signal WR_MA                : std_logic;
    signal RD_MA                : std_logic;

    -- DTU MA Stage (DFFs -> DTU)
    signal DBInMode_WB          : integer range DBINMODE_CNT-1 downto 0;
    signal DataAccessMode_WB    : integer range DATAACCESSMODE_CNT-1 downto 0;
    signal WR_WB                : std_logic;
    signal RD_WB                : std_logic;

    ---------------------------------------------------------------------------
    -- CU Signals
    ---------------------------------------------------------------------------

    -- Pipeline some bits of IR to use as offset to ALU, PAU, DAU
    signal IR_ID : std_logic_vector(INST_SIZE-1 downto 0);
    signal IR_EX : std_logic_vector(11 downto 0);   -- max offset is only 12-bits
    signal IR_MA : std_logic_vector(11 downto 0);   

    -- Pipeline when to update IR (fed back into CU)
    signal UpdateIR_ID : std_logic;
    signal UpdateIR_EX : std_logic;
    signal UpdateIR_MA : std_logic;
    signal UpdateIR_WB : std_logic;

    -- Pipeline when to update SR (fed back into CU)
    signal UpdateSR_ID : std_logic;
    signal UpdateSR_EX : std_logic;
    signal UpdateSR_MA : std_logic;
    signal UpdateSR_WB : std_logic;
    signal SRSel_ID    : integer range SRSEL_CNT-1 downto 0;
    signal SRSel_EX    : integer range SRSEL_CNT-1 downto 0;
    signal SRSel_MA    : integer range SRSEL_CNT-1 downto 0;
    signal SRSel_WB    : integer range SRSEL_CNT-1 downto 0;

    -- Pipeline read-modify-write (RMW) command
    signal RMW_ID : std_logic;
    signal RMW_EX : std_logic;
    signal RMW_MA : std_logic;
    signal RMW_WB : std_logic;

    -- Non-pipelined outputs
    signal SR : std_logic_vector(REG_SIZE-1 downto 0);
    signal TempReg : std_logic_vector(31 downto 0);
    signal TempReg2 : std_logic_vector(31 downto 0);

    ---------------------------------------------------------------------------
    -- Top-Level Control Signals
    ---------------------------------------------------------------------------

    -- Pipeline data bus output control signals to determine source of DBOut
    signal DBOutSel_ID : integer range DBOUTSEL_CNT-1 downto 0;
    signal DBOutSel_EX : integer range DBOUTSEL_CNT-1 downto 0;
    signal DBOutSel_MA : integer range DBOUTSEL_CNT-1 downto 0;
    signal DBOutSel_WB : integer range DBOUTSEL_CNT-1 downto 0;

    -- Pipeline address bus output control signals to determine source of AB
    signal ABOutSel_ID : integer range 1 downto 0;
    signal ABOutSel_EX : integer range 1 downto 0;
    signal ABOutSel_MA : integer range 1 downto 0;
    signal ABOutSel_WB : integer range 1 downto 0;

    -- Create muxes for data forwarding to avoid data bus and address bus contentions
    signal DBMux : std_logic_vector(DATA_BUS_SIZE-1 downto 0); -- select DB or delayed DB
    signal ABMux : std_logic_vector(1 downto 0);               -- select AB or delayed AB

    -- Create 1 clock delays for data bus and address bus (useful for data forwarding)
    signal DB_Delayed : std_logic_vector(DATA_BUS_SIZE-1 downto 0);  -- delayed DB by 1 clock
    signal AB_Delayed : std_logic_vector(1 downto 0);                -- delayed AB by 1 clock

    -- Pipeline branch type selection so addresses are calculated in EX stage
    signal BranchSel_ID : integer range BRANCHSEL_CNT-1 downto 0;
    signal BranchSel_EX : integer range BRANCHSEL_CNT-1 downto 0;

    -- Create muxes to select source and offset to PAU (needed for branch control hazards)
    signal PAU_SrcSel_Mux       : integer range PAU_SRC_CNT - 1 downto 0;
    signal PAU_OffsetSel_Mux    : integer range PAU_OFFSET_CNT - 1 downto 0;
    signal PAU_UpdatePC_Mux     : std_logic;

    -- Create mux to select when registers should be written to
    signal RegStore_Mux     : std_logic;
    signal RegAxStore_Mux   : std_logic;

    -- Mux to determine which source to use to update instruction register (IR)
    signal UpdateIR_Mux : std_logic;

    -- Pipeline signal that indicates when write back state should be used
    signal UseWB_ID : std_logic;
    signal UseWB_EX : std_logic;
    signal UseWB_MA : std_logic;
    signal UseWB_WB : std_logic;

    -- Data bus inputs and outputs
    signal DBIn     : std_logic_vector(DATA_BUS_SIZE-1 downto 0);
    signal DBOut    : std_logic_vector(DATA_BUS_SIZE-1 downto 0);

    -- Indicate when a branch should be taken
    signal TakeBranch : std_logic;

    -- Indicate when stages of pipeline should be stalled
    signal StallPL_ID : std_logic;
    signal StallPL_EX : std_logic;
    signal StallPL_MA : std_logic;
    signal StallPL_WB : std_logic;

    -- Indicate when the pipeline should be flushed
    signal FlushPL : std_logic;

begin

    -- Select address to be either address output by PAU or DAU
    AB <= PAU_ProgAddr when ABOutSel_MA = ABOutSel_Prog else
          DAU_DataAddr when ABOutSel_MA = ABOutSel_Data else
          (others => 'X');

    -- Select data to output to data bus
    DBOut <= ALU_Result when DBOutSel_MA = DBOutSel_Result else
             GBR        when DBOutSel_MA = DBOutSel_GBR    else
             VBR        when DBOutSel_MA = DBOutSel_VBR    else
             SR         when DBOutSel_MA = DBOutSel_SR     else
             PR         when DBOutSel_MA = DBOutSel_PR     else
             PC_ID      when DBOutSel_MA = DBOutSel_PC     else
             (others => 'X');

    -- Update the CU data bus input either normal or memory access stalled input
    DBMux <= DB_Delayed when UpdateIR_MA = '0' and UpdateSR_EX = '0' else DB;
    ABMux <= AB_Delayed when UpdateIR_MA = '0' else AB(1 downto 0);

    -- These muxes prevent registers from storing values on multiple clocks
    RegStore_Mux <= RegStore_EX when UseWB_WB = '0' else RegStore_WB;
    RegAxStore_Mux <= RegAxStore_MA when UseWB_WB = '0' else RegAxStore_WB;


    UpdateIR_Mux <= UpdateIR_EX;

    -- Combinational logic to handle branching and control hazards
    Branching  : process (all)
    begin

        -- Check if branch should be taken
        if BranchSel_EX = BranchSel_BF or BranchSel_EX = BranchSel_BFS then
            TakeBranch <= '1' when SR(0) = '0' else '0';    -- Branch when T-bit clear
        elsif BranchSel_EX = BranchSel_BT or BranchSel_EX = BranchSel_BTS then
            TakeBranch <= '1' when SR(0) = '1' else '0';    -- Branch when T-bit set
        elsif BranchSel_EX /= BranchSel_None then
            TakeBranch <= '1';  -- Always branch
        else
            TakeBranch <= '0';  -- Not a branch instruction so don't branch
        end if;

        -- Flush pipeline if branching without a slot instruction
        FlushPL <= '1' when TakeBranch = '1' and (BranchSel_EX = BranchSel_BF or BranchSel_EX = BranchSel_BT) else '0';

        -- Select PAU source to calculate address to branch to (if branching)
        if TakeBranch = '1' then
            if (BranchSel_EX = BranchSel_Direct) then
                PAU_SrcSel_Mux <= PAU_AddrPC_EX;    -- pipelined PC value
            elsif (BranchSel_EX = BranchSel_RET) then
                PAU_SrcSel_Mux <= PAU_AddrPR;       -- PR
            elsif (BranchSel_EX = BranchSel_Indirect) then
                PAU_SrcSel_Mux <= PAU_AddrZero;     -- zero since address in offset reg
            else
                PAU_SrcSel_Mux <= PAU_AddrPC_EX;    -- pipelined PC value
            end if;
        else
            PAU_SrcSel_Mux <= PAU_SrcSel_EX;        -- normal PC offset
        end if;

        -- Mux to select PAU offset to calculate address to branch to if branching
        PAU_OffsetSel_Mux <= PAU_OffsetSel_EX when TakeBranch = '1' and BranchSel_EX /= BranchSel_None else
                             PAU_OffsetWord;

        PAU_UpdatePC_Mux <= PAU_UpdatePC_EX;

    end process;


    -- Insert DFFs into pipeline and give default values upon reset or pipeline flush
    Pipeline : process (clock)
    begin
        -- Pass on instructions from one stage to the stage
        if rising_edge(clock) then
        
            -- Define initial values upon reset
            if reset = '0' then

                -- Set pipeline values to read in first instruction
                -- Essentially fill pipeline with NOP control signals

                -- EX stage
                DBInMode_EX <= DBInMode_Unsigned;
                DataAccessMode_EX <= DataAccessMode_WORD;
                WR_EX <= '1';
                RD_EX <= '0';
                UpdateIR_EX <= '1';
                UpdateIR_MA <= '1';
                ABOutSel_EX <= ABOutSel_Prog;
                
                -- MA stage
                DBInMode_MA <= DBInMode_Unsigned;
                DataAccessMode_MA <= DataAccessMode_WORD;
                WR_MA <= '1';
                RD_MA <= '0';
                ABOutSel_MA <= ABOutSel_Prog;
        
            else
                    
                ---------------------------------------------------------------
                -- ID to EX DFFs
                ---------------------------------------------------------------

                -- Pipelined signals that cannot be stalled. Some are given
                -- default values for when pipeline is flushed.
                -- Avoid contentions on address bus when there is a memory access
                -- before/after the branch instruction
                if (TakeBranch = '1' and ABOutSel_MA = ABOutSel_Data) then
                    BranchSel_EX <= BranchSel_EX;
                    PAU_OffsetSel_EX <= PAU_OffsetSel_ID;
                else
                    BranchSel_EX <= BranchSel_ID when FlushPL = '0' else BranchSel_None;
                    PAU_OffsetSel_EX    <= PAU_OffsetSel_ID when TakeBranch = '0' else PAU_OffsetWord; 
                end if;

                                    -- PAU signals
                    PAU_UpdatePC_EX     <= PAU_UpdatePC_ID;
                    PAU_PRSel_EX        <= PAU_PRSel_ID when FlushPL = '0' else PRSel_None;
                    PAU_IncDecSel_EX    <= PAU_IncDecSel_ID;
                    PAU_IncDecBit_EX    <= PAU_IncDecBit_ID;
                    PAU_PrePostSel_EX   <= PAU_PrePostSel_ID;
                    PC_EX               <= PC_ID when FlushPL = '0' else AB;
                    PAU_SrcSel_EX       <= PAU_SrcSel_ID when TakeBranch = '0' else PAU_AddrPC;

  
                StallPL_EX <= StallPL_ID;

                -- DTU signals
                DBInMode_EX <= DBInMode_ID;
                DataAccessMode_EX <= DataAccessMode_ID;
                WR_EX <= WR_ID when FlushPL = '0' else '1';
                RD_EX <= RD_ID when FlushPL = '0' else '0';

                -- CU signals
                UpdateIR_EX         <= UpdateIR_ID when FlushPL = '0' else '1';

                -- Top-level signals
                DBOutSel_EX         <= DBOutSel_ID;
                ABOutSel_EX         <= ABOutSel_ID;
                UseWB_EX            <= UseWB_ID;
                RMW_EX              <= RMW_ID;

                -- Stall some signals when neccessary. Some are given default
                -- values for when pipeline is flushed.
                if StallPL_EX = '0' then

                    -- ALU signals
                    ALUOpASel_EX    <= ALUOpASel_ID;
                    ALUOpBSel_EX    <= ALUOpBSel_ID;
                    ALU_FCmd_EX     <= ALU_FCmd_ID;
                    ALU_CinCmd_EX   <= ALU_CinCmd_ID;
                    ALU_SCmd_EX     <= ALU_SCmd_ID;
                    ALU_ALUCmd_EX   <= ALU_ALUCmd_ID;
                    ALU_TbitOp_EX   <= ALU_TbitOp_ID;

                    -- RegArray signals
                    RegInSel_EX         <= RegInSel_ID;
                    RegStore_EX         <= RegStore_ID when FlushPL = '0' else '0';
                    RegASel_EX          <= RegASel_ID;
                    RegBSel_EX          <= RegBSel_ID;
                    RegAxInSel_EX       <= RegAxInSel_ID;
                    RegAxInDataSel_EX   <= RegAxInDataSel_ID;
                    RegAxStore_EX       <= RegAxStore_ID when FlushPL = '0' else '0';
                    RegA1Sel_EX         <= RegA1Sel_ID;
                    RegOpSel_EX         <= RegOpSel_ID;

                    -- DAU signals
                    DAU_SrcSel_EX       <= DAU_SrcSel_ID when FlushPL = '0' else DAU_SrcSel_EX;
                    DAU_OffsetSel_EX    <= DAU_OffsetSel_ID when FlushPL = '0' else DAU_OffsetSel_EX;                    
                    DAU_Offset4_EX      <= DAU_Offset4_ID when FlushPL = '0' else DAU_Offset4_EX;
                    DAU_Offset8_EX      <= DAU_Offset8_ID when FlushPL = '0' else DAU_Offset8_EX;                    
                    DAU_IncDecSel_EX    <= DAU_IncDecSel_ID when FlushPL = '0' else DAU_IncDecSel_EX;
                    DAU_IncDecBit_EX    <= DAU_IncDecBit_ID when FlushPL = '0' else DAU_IncDecBit_EX;
                    DAU_PrePostSel_EX   <= DAU_PrePostSel_ID when FlushPL = '0' else DAU_PrePostSel_EX;
                    DAU_GBRSel_EX       <= DAU_GBRSel_ID when FlushPL = '0' else GBRSel_None;
                    DAU_VBRSel_EX       <= DAU_VBRSel_ID when FlushPL = '0' else VBRSel_None;

                    -- CU signals
                    UpdateSR_EX <= UpdateSR_ID when FlushPL = '0' else '0';
                    SRSel_EX    <= SRSel_ID;

                    -- Top-level signals
                    IR_EX   <= IR_ID(11 downto 0);

                end if;

                ---------------------------------------------------------------
                -- EX to MA DFFs
                ---------------------------------------------------------------

                -- Pipelined signals that cannot be stalled. Some are given
                -- default values for when pipeline is flushed.

                -- Instruction register data
                IR_MA <= IR_EX(11 downto 0);

                -- DAU control signals
                DAU_SrcSel_MA       <= DAU_SrcSel_EX;
                DAU_OffsetSel_MA    <= DAU_OffsetSel_EX;
                DAU_Offset4_MA      <= DAU_Offset4_EX;
                DAU_Offset8_MA      <= DAU_Offset8_EX;
                DAU_IncDecSel_MA    <= DAU_IncDecSel_EX;
                DAU_IncDecBit_MA    <= DAU_IncDecBit_EX;
                DAU_PrePostSel_MA   <= DAU_PrePostSel_EX;
                DAU_GBRSel_MA       <= DAU_GBRSel_EX;
                DAU_VBRSel_MA       <= DAU_VBRSel_EX;

                -- Top-level signals
                DB_Delayed  <= DB;
                AB_Delayed  <= AB(1 downto 0);

                    -- DTU signals
                DBInMode_MA         <= DBInMode_EX;
                DataAccessMode_MA   <= DataAccessMode_EX;
                WR_MA               <= WR_EX;
                RD_MA               <= RD_EX;

                -- CU signals
                UpdateIR_MA <= UpdateIR_EX when FlushPL = '0' else '1';

                -- Top-level signals
                DBOutSel_MA     <= DBOutSel_EX;
                ABOutSel_MA     <= ABOutSel_EX;
                UseWB_MA        <= UseWB_EX;
                RMW_MA          <= RMW_EX;

                StallPL_MA <= StallPL_EX;

                ---------------------------------------------------------------
                -- MA to WB DFFs
                ---------------------------------------------------------------
                UseWB_WB    <= UseWB_MA;
                RMW_WB      <= RMW_MA;

                StallPL_WB <= StallPL_MA;

            end if;

        end if;

    end process;


-- SH2 CPU Component Implementation and Port Mapping
--  Create the all SH2 CPU component and map the ports to the internal signals.

    -- Create 32-bit ALU for standard logic and arithmetic operations
    SH2_ALU : ALU
        port map (
            -- Operand signals (inputs)
            RegA        => RegA,
            RegB        => RegB,
            TempReg     => TempReg2,
            Imm         => IR_EX(7 downto 0),
            DBIn        => DBIn,
            SR0         => SR(0),

            -- Control signals (inputs)
            ALUOpASel   => ALUOpASel_EX,
            ALUOpBSel   => ALUOpBSel_EX,
            FCmd        => ALU_FCmd_EX,
            CinCmd      => ALU_CinCmd_EX,
            SCmd        => ALU_SCmd_EX,
            ALUCmd      => ALU_ALUCmd_EX,

            -- Output signals            
            TbitOp      => ALU_TbitOp_EX,
            Result      => ALU_Result,
            Tbit        => ALU_Tbit
        );

    -- Create 32-bit register array with general purpose registers R0-R15
    SH2_RegArray : RegArray
        port map (
            -- RegIn input
            Result          => ALU_Result,

            -- RegAxIn inputs
            DataAddrID      => DAU_AddrIDOut,
            DataAddr        => DAU_DataAddr,
            SR              => SR,
            GBR             => GBR,
            VBR             => VBR,
            PR              => PR,

            -- Control signals (inputs)
            RegInSel        => RegInSel_EX,
            RegStore        => RegStore_Mux,
            RegASel         => RegASel_EX,
            RegBSel         => RegBSel_EX,
            RegAxInSel      => RegAxInSel_EX,
            RegAxInDataSel  => RegAxInDataSel_EX,
            RegAxStore      => RegAxStore_Mux,
            RegA1Sel        => RegA1Sel_EX,
            RegOpSel        => RegOpSel_EX,
            CLK             => clock,

            -- Register outputs
            RegA            => RegA,
            RegB            => RegB,
            RegA1           => RegA1
        );

    -- Create Program Memory Access Unit (PAU)
    SH2_PAU : PAU
        port map (
            -- Control signals
            SrcSel     => PAU_SrcSel_Mux,
            OffsetSel  => PAU_OffsetSel_Mux,
            UpdatePC   => PAU_UpdatePC_Mux,
            PRSel      => PAU_PRSel_EX,
            IncDecSel  => PAU_IncDecSel_EX,
            IncDecBit  => PAU_IncDecBit_EX,
            PrePostSel => PAU_PrePostSel_EX,

            -- Source inputs
            DB         => DB,
            PC_EX      => PC_EX,

            -- Offset inputs
            Offset8    => IR_EX(7 downto 0),
            Offset12   => IR_EX(11 downto 0),
            OffsetReg  => RegA1,
            TempReg    => TempReg,

            -- System signal
            CLK        => clock,
            RESET      => reset,

            -- Output signals
            ProgAddr   => PAU_ProgAddr,
            PC         => PC_ID,
            PR         => PR
        );

    -- Create Data Memory Access Unit (DAU)
    SH2_DAU : DAU
        port map (
            -- Source inputs
            PC         => PC_ID,
            Rn         => RegA1,

            -- Offset inputs
            Offset4    => IR_EX(3 downto 0),
            Offset8    => IR_EX(7 downto 0),
            R0         => RegA,

            -- Data inputs
            DB         => DB,

            -- Control signals
            SrcSel     => DAU_SrcSel_EX,
            OffsetSel  => DAU_OffsetSel_EX,
            IncDecSel  => DAU_IncDecSel_EX,
            IncDecBit  => DAU_IncDecBit_EX,
            PrePostSel => DAU_PrePostSel_EX,
            GBRSel     => DAU_GBRSel_EX,
            VBRSel     => DAU_VBRSel_EX,
            CLK        => clock,
            RST        => Reset,

            -- Output signals
            AddrIDOut  => DAU_AddrIDOut,
            DataAddr   => DAU_DataAddr,
            GBR        => GBR,
            VBR        => VBR
        );

    -- Create Data Transfer Unit (DTU) to interface with memory
    SH2_DTU : DTU
        port map (
            -- Data input
            DBOut           => DBOut,

            -- Control inputs
            AB              => AB(1 downto 0),
            RD              => RD_MA,
            WR              => WR_MA,
            DataAccessMode  => DataAccessMode_MA,
            DBInMode        => DBInMode_MA,
            CLK             => clock,

            -- Control outputs
            DBIn            => DBIn,
            WE0             => WE0,
            WE1             => WE1,
            WE2             => WE2,
            WE3             => WE3,
            RE0             => RE0,
            RE1             => RE1,
            RE2             => RE2,
            RE3             => RE3,

            -- In/Out data bus
            DB              => DB
        );

    -- Control Unit (CU)
    SH2_CU : CU
        port map (
            
            -- CU Input Signals
            CLK         => clock,
            RST         => reset,
            DB          => DBMux,
            AB          => ABMux,
            RegB        => RegB,
            Result      => ALU_Result,

            -- CU Registers
            SR          => SR,
            IR          => IR_ID,
            Tbit        => ALU_Tbit,
            TempReg     => TempReg,
            TempReg2    => TempReg2,

            -- CU Output Signals
            UpdateIR   => UpdateIR_ID,
            UpdateSR   => UpdateSR_ID,
            SRSel      => SRSel_ID,
            SRSel_EX   => SRSel_EX,

            -- ALU Signals
            ALUOpASel   => ALUOpASel_ID,
            ALUOpBSel   => ALUOpBSel_ID,
            FCmd        => ALU_FCmd_ID,
            CinCmd      => ALU_CinCmd_ID,
            SCmd        => ALU_SCmd_ID,
            ALUCmd      => ALU_ALUCmd_ID,
            TbitOp      => ALU_TbitOp_ID,

            -- PAU Signals
            PAU_SrcSel      => PAU_SrcSel_ID,
            PAU_OffsetSel   => PAU_OffsetSel_ID,
            PAU_UpdatePC    => PAU_UpdatePC_ID,
            PAU_PRSel       => PAU_PRSel_ID,
            PAU_IncDecSel   => PAU_IncDecSel_ID,
            PAU_IncDecBit   => PAU_IncDecBit_ID,
            PAU_PrePostSel  => PAU_PrePostSel_ID,

            -- DAU Signals
            DAU_SrcSel      => DAU_SrcSel_ID,
            DAU_OffsetSel   => DAU_OffsetSel_ID,
            DAU_IncDecSel   => DAU_IncDecSel_ID,
            DAU_IncDecBit   => DAU_IncDecBit_ID,
            DAU_PrePostSel  => DAU_PrePostSel_ID,
            DAU_GBRSel      => DAU_GBRSel_ID,
            DAU_VBRSel      => DAU_VBRSel_ID,

            -- RegArray Signals
            RegInSel        => RegInSel_ID,
            RegStore        => RegStore_ID,
            RegASel         => RegASel_ID,
            RegBSel         => RegBSel_ID,
            RegAxInSel      => RegAxInSel_ID,
            RegAxInDataSel  => RegAxInDataSel_ID,
            RegAxStore      => RegAxStore_ID,
            RegA1Sel        => RegA1Sel_ID,
            RegOpSel        => RegOpSel_ID,

            -- DTU signals
            RD => RD_ID,
            WR => WR_ID,
            DataAccessMode => DataAccessMode_ID,
            DBInMode => DBInMode_ID,

            -- IO signals
            DBOutSel    => DBOutSel_ID,
            ABOutSel    => ABOutSel_ID,

            -- Pipeline signals
            StallPL => StallPL_ID,
            UpdateIR_EX => UpdateIR_Mux,
            UpdateSR_EX => UpdateSR_EX,
            TakeBranch => TakeBranch,
            RMW => RMW_ID,
            UseWB => UseWB_ID,
            BranchSel => BranchSel_ID
        );

end structural;