----------------------------------------------------------------------------
--
--  SH-2 Control Unit
--
--  This file contains the control unit (CU) implementation for a SH-2 processor.
--  It decodes instructions and generates control signals for the ALU, PAU, DAU,
--  RegArray, DTU, and top-level muxes. It also includes a FSM for instruction
--  sequencing and control
--
--  Packages included are:
--   CUConstants - constants for control signal values
--
--  Entities included are:
--   CU - control unit    
--
--  Revision History:
--     18 April 2025    Garrett Knuf    Initial revision.
--     20 April 2025    Garrett Knuf    Add autogen markers for instruction decoding.
--     24 April 2025    Garrett Knuf    Add FSM.
--     12 May 2025      Garrett Knuf    Fix bugs in decoding.
--     15 May 2025      Garrett Knuf    Optimize logic.
--
----------------------------------------------------------------------------

--
-- Package containing constants for the control unit.
--

library ieee;
use ieee.std_logic_1164.all;
use work.GenericConstants.all;
use work.RegArrayConstants.all;

package CUConstants is

    -- RegInSel - select where to save input to RegIn
    constant REGINSELCMD_CNT   : integer := 3;
    constant RegInSelCmd_Rn    : integer range REGINSELCMD_CNT-1 downto 0 := 0;    -- generic register
    constant RegInSelCmd_R0    : integer range REGINSELCMD_CNT-1 downto 0 := 1;    -- register R0
    constant RegInSelCmd_R15   : integer range REGINSELCMD_CNT-1 downto 0 := 2;    -- register R15

    -- RegASelCmd - select what RegA outputs
    constant RegASelCmd_Rn : integer range 2 downto 0 := 0;     -- generic register
    constant RegASelCmd_DB : integer range 2 downto 0 := 1;     -- databus
    constant RegASelCmd_R0 : integer range 2 downto 0 := 2;     -- register R0

    -- RegBSelCmd - select what RegB outputs
    constant RegBSelCmd_Rm : integer range 2 downto 0 := 0;     -- generic register
    constant RegBSelCmd_R0 : integer range 2 downto 0 := 1;     -- register R0
    constant RegBSelCmd_Rn : integer range 2 downto 0 := 2;     -- generic register
    
    -- RegA1SelCmd - select what RegA1 outputs
    constant RegA1SelCmd_CNT : integer := 4;
    constant RegA1SelCmd_Rn  : integer range RegA1SelCmd_CNT-1 downto 0 := 0;   -- generic register
    constant RegA1SelCmd_Rm  : integer range RegA1SelCmd_CNT-1 downto 0 := 1;   -- generic register
    constant RegA1SelCmd_R0  : integer range RegA1SelCmd_CNT-1 downto 0 := 2;   -- R0
    constant RegA1SelCmd_R15 : integer range RegA1SelCmd_CNT-1 downto 0 := 3;   -- R15

    -- RegAxInSelCmd - select what RegA1 outputs
    constant RegAxInSelCmd_CNT : integer := 4;
    constant RegAxInSelCmd_Rn  : integer range RegAxInSelCmd_CNT-1 downto 0 := 0;   -- generic register
    constant RegAxInSelCmd_Rm  : integer range RegAxInSelCmd_CNT-1 downto 0 := 1;   -- generic register
    constant RegAxInSelCmd_R0  : integer range RegAxInSelCmd_CNT-1 downto 0 := 2;   -- R0
    constant RegAxInSelCmd_R15 : integer range RegAxInSelCmd_CNT-1 downto 0 := 3;   -- R15

    -- DBOutSel - select output of databus
    constant DBOUTSEL_CNT    : integer := 6;
    constant DBOutSel_Result : integer range DBOUTSEL_CNT-1 downto 0 := 0;  -- ALU result
    constant DBOutSel_SR     : integer range DBOUTSEL_CNT-1 downto 0 := 1;  -- status reg
    constant DBOutSel_GBR    : integer range DBOUTSEL_CNT-1 downto 0 := 2;  -- GBR
    constant DBOutSel_VBR    : integer range DBOUTSEL_CNT-1 downto 0 := 3;  -- VBR
    constant DBOutSel_PR     : integer range DBOUTSEL_CNT-1 downto 0 := 4;  -- PR
    constant DBOutSel_PC     : integer range DBOUTSEL_CNT-1 downto 0 := 5;  -- PC

    -- ABSel - select output of address bus
    constant ABOutSel_Prog : integer range 1 downto 0 := 0; -- PAU address
    constant ABOutSel_Data : integer range 1 downto 0 := 1; -- DAU address

    -- TempRegSel - select value to put into temporary register
    constant TempRegSel_CNT      : integer := 5;
    constant TempRegSel_Offset8  : integer range TempRegSel_CNT-1 downto 0 := 0;
    constant TempRegSel_Offset12 : integer range TempRegSel_CNT-1 downto 0 := 1;
    constant TempRegSel_RegB     : integer range TempRegSel_CNT-1 downto 0 := 2;
    constant TempRegSel_Result   : integer range TempRegSel_CNT-1 downto 0 := 3;
    constant TempRegSel_DataBus  : integer range TempRegSel_CNT-1 downto 0 := 4;

    -- TempReg2Sel - select value to put into temporary register 2
    constant TempReg2Sel_CNT      : integer := 2;
    constant TempReg2Sel_Result   : integer range TempRegSel_CNT-1 downto 0 := 0;
    constant TempReg2Sel_DB       : integer range TempRegSel_CNT-1 downto 0 := 1;

    -- Bit indices of SR
    constant StatusReg_Tbit     : integer := 0; -- T bit
    constant StatusReg_Sbit     : integer := 1; -- S bit
    constant StatusReg_I0bit    : integer := 4; -- Interrupt mask I0
    constant StatusReg_I1bit    : integer := 5; -- Interrupt mask I1
    constant StatusReg_I2bit    : integer := 6; -- Interrupt mask I2
    constant StatusReg_I3bit    : integer := 7; -- Interrupt mask I3
    constant StatusReg_Qbit     : integer := 8; -- Q bit
    constant StatusReg_Mbit     : integer := 9; -- M bit

    -- SRSel - select value to load into SR
    constant SRSEL_CNT  : integer := 4;
    constant SRSel_Tbit : integer range SRSEL_CNT-1 downto 0 := 0;  -- Set Tbit
    constant SRSel_DB   : integer range SRSEL_CNT-1 downto 0 := 1;  -- Set to DB
    constant SRSel_Reg  : integer range SRSEL_CNT-1 downto 0 := 2;  -- Set to register
    constant SRSel_Tmp2 : integer range SRSEL_CNT-1 downto 0 := 3;  -- Set to temporary reg 2

    constant unused : integer := 0;

end package;


--
-- This architecture implements the finite state machine (FSM) and instruction
-- decoding logic for the SH-2 control unit. It generates approprate
-- control signals for:
--  ALU operation selection and operand routing
--  Program address updates via the PAU
--  Data addres updates via the DAU
--  Register access and storage
--  Memory and I/O control
--  Special handling for T-bit and SR register operations
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.GenericConstants.all;
use work.DTUConstants.all;
use work.CUConstants.all;
use work.ALUConstants.all;
use work.GenericALUConstants.all;
use work.MemUnitConstants.all;
use work.DAUConstants.all;
use work.PAUConstants.all;
use work.RegArrayConstants.all;
use work.OpcodeConstants.all;

entity CU is

    port (
     -- CU Input Signals
        CLK     : in    std_logic;                                      -- system clock
        RST     : in    std_logic;                                      -- system reset
        DB      : in    std_logic_vector(DATA_BUS_SIZE - 1 downto 0);   -- data bus
        AB      : in    std_logic_vector(1 downto 0);                   -- address bus (least 2 significant bits)
        Result  : in    std_logic_vector(LONG_SIZE - 1 downto 0);       -- ALU result
        Tbit    : in    std_logic;                                      -- Tbit from ALU
        RegB    : in    std_logic_vector(REG_SIZE - 1 downto 0);

        -- CU Registers
        IR      : out   std_logic_vector(INST_SIZE - 1 downto 0) := x"DEAD";    -- instruction register
        SR      : out std_logic_vector(REG_SIZE - 1 downto 0);                  -- status register
        TempReg : out std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);             -- temporary register
        TempReg2 : out std_logic_vector(ADDR_BUS_SIZE - 1 downto 0);            -- secondary temp register
        
        -- CU Output Signals
        UpdateIR  : out   std_logic;    -- update instruction register (used to delay pipeline during data access)
        UpdateSR  : out   std_logic;

        -- ALU Control Signals
        ALUOpASel   : out     integer range ALUOPASEL_CNT-1 downto 0 := 0;  -- select operand A
        ALUOpBSel   : out     integer range ALUOPBSEL_CNT-1 downto 0 := 0;  -- select operand B
        FCmd        : out     std_logic_vector(3 downto 0);                 -- Fblock control
        CinCmd      : out     std_logic_vector(1 downto 0);                 -- carry in
        SCmd        : out     std_logic_vector(2 downto 0);                 -- shift block control
        ALUCmd      : out     std_logic_vector(1 downto 0);                 -- output mux
        TbitOp      : out     std_logic_vector(3 downto 0);                 -- tbit control

        -- PAU Control Signals
        PAU_SrcSel      : out   integer range PAU_SRC_CNT - 1 downto 0;     -- select address source
        PAU_OffsetSel   : out   integer range PAU_OFFSET_CNT - 1 downto 0;  -- select offset source
        PAU_UpdatePC    : out   std_logic;                                  -- update PC
        PAU_PRSel       : out   integer range PRSEL_CNT-1 downto 0;         -- select PR control
        PAU_IncDecSel   : out   std_logic;                                  -- select inc/dec
        PAU_IncDecBit   : out   integer range 2 downto 0;                   -- select inc/dec bit
        PAU_PrePostSel  : out   std_logic;                                  -- select pre/post

        -- DAU Control Signals
        DAU_SrcSel      : out   integer range DAU_SRC_CNT - 1 downto 0;     -- select address source
        DAU_OffsetSel   : out   integer range DAU_OFFSET_CNT - 1 downto 0;  -- select offset source
        DAU_IncDecSel   : out   std_logic;                                  -- select inc/dec
        DAU_IncDecBit   : out   integer range 2 downto 0;                   -- select inc/dec bit
        DAU_PrePostSel  : out   std_logic;                                  -- select pre/post
        DAU_GBRSel      : out   integer range GBRSEL_CNT-1 downto 0;        -- select GBR load
        DAU_VBRSel      : out   integer range VBRSEL_CNT-1 downto 0;        -- select VBR load

        -- RegArray Control Signals
        RegInSel        : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select input reg
        RegStore        : out   std_logic;                                      -- store input reg
        RegASel         : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select output RegA
        RegBSel         : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select output regB
        RegAxInSel      : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select address input reg
        RegAxInDataSel  : out   integer range REGAXINDATASEL_CNT - 1 downto 0;  -- select data to address input
        RegAxStore      : out   std_logic;                                      -- store address input
        RegA1Sel        : out   integer  range REGARRAY_RegCnt - 1 downto 0;    -- select address reg output
        RegOpSel        : out   integer  range REGOPSEL_CNT - 1 downto 0;       -- select special reg operation
    
        -- IO Control signals
        DBOutSel : out integer range DBOUTSEL_CNT-1 downto 0;   -- select databus output
        ABOutSel : out integer range 1 downto 0;                -- select addressbus output
        DBInMode : out integer range 1 downto 0;                -- select sign/unsigned databus read
        RD     : out   std_logic;                               -- read (active-low)
        WR     : out   std_logic;                               -- write (active-low)
        DataAccessMode : out integer range 2 downto 0;          -- align bytes, words, long

        -- Pipeline control signals
        UpdateIR_EX : in std_logic;    -- pipelined signal to update IR
        UpdateSR_EX : in std_logic;    -- pipelined control signal to update SR or not
        ForceNormalStateNext : in std_logic
    );


end CU;

architecture behavioral of CU is

    -- Finite-state machine (FSM) states
    constant Normal             : integer := 0; -- fetch next instruction while executing current
    constant WaitForFetch       : integer := 1; -- one clock wait to fetch next instruction
    constant BranchSlot         : integer := 2; -- branch slot to reg+offset
    constant BranchSlotRet      : integer := 3; -- branch slot when returning from function call
    constant BranchSlotDirect   : integer := 4; -- branch slot to offset
    constant BootReadSP         : integer := 5; -- read stack pointer from vec table on boot
    constant BootWaitForFetch   : integer := 6; -- fetch first instruction to run after boot sequence
    constant WriteBack          : integer := 7; -- write a value from temp reg back to memory
    constant TRAPA_PushPC       : integer := 8; -- push PC onto stack
    constant TRAPA_ReadVector   : integer := 9; -- read vector address
    constant RTE_PopSR          : integer := 10; -- pop SR from stack
    constant RTE_Slot           : integer := 11; -- RTE branch slot
    constant Sleep              : integer := 12; -- idle (no code executing)
    constant STATE_CNT          : integer := 13; -- total number of states

    signal NextState : integer range STATE_CNT-1 downto 0;      -- state to transition to on next clock
    signal CurrentState : integer range STATE_CNT-1 downto 0;   -- current state being executed

    -- CU internal control signals
    signal SRSel : integer range SRSEL_CNT-1 downto 0;                  -- select input to status register

    signal RegInSelCmd : integer range REGARRAY_RegCnt-1 downto 0;      -- select register for RegArray input
    signal RegASelCmd : integer range REGARRAY_RegCnt-1 downto 0;       -- select register for RegArray RegA
    signal RegBSelCmd : integer range REGARRAY_RegCnt-1 downto 0;       -- select register for RegArray RegB
    signal RegAxInSelCmd : integer range REGARRAY_RegCnt-1 downto 0;    -- select register for RegArray address input 
    signal RegA1SelCmd : integer range REGARRAY_RegCnt-1 downto 0;      -- select register for RegArray RegA1

    signal UpdateTempReg : std_logic;                                   -- control signal to update TempReg or not
    signal TempRegSel : integer range TempRegSel_CNT-1 downto 0;        -- select temporary register input
    signal TempRegMuxOut : std_logic_vector(REG_SIZE-1 downto 0);       -- mux input to TempReg
    signal TempReg2MuxOut : std_logic_vector(REG_SIZE-1 downto 0);      -- mux input to TempReg2
    signal UpdateTempReg2 : std_logic;                                  -- update secondary temporary register
    signal TempReg2Sel  : integer range TempReg2Sel_CNT-1 downto 0;     -- secondary temporary register select
    
begin

    -- Signal to set temporary register 1 to
    TempRegMuxOut <= (31 downto 9 => IR(7)) & IR(7 downto 0) & '0' when TempRegSel = TempRegSel_Offset8 else
                     (31 downto 13 => IR(11)) & IR(11 downto 0) & '0' when TempRegSel = TempRegSel_Offset12 else
                     RegB when TempRegSel = TempRegSel_RegB else
                     Result when TempRegSel = TempRegSel_Result else
                     DB when TempRegSel = TempRegSel_DataBus else
                     (others => 'X');

    -- Signal to set temporary register 2 to
    TempReg2MuxOut <= DB     when TempReg2Sel = TempReg2Sel_DB else
                      Result when TempReg2Sel = TempReg2Sel_Result else
                      (others => 'X');

    -- Select registers to access in register array
    RegInSel <= to_integer(unsigned(IR(11 downto 8)))   when RegInSelCmd = RegInSelCmd_Rn else
                R15                                     when RegInSelCmd = RegInSelCmd_R15 else
                R0;

    RegASel <= to_integer(unsigned(IR(11 downto 8)))    when RegASelCmd = RegASelCmd_Rn else R0;

    RegBSel <= to_integer(unsigned(IR(7 downto 4)))     when RegBSelCmd = RegBSelCmd_Rm else
               to_integer(unsigned(IR(11 downto 8)))    when RegBSelCmd = RegBSelCmd_Rn else R0;

    RegA1Sel <= to_integer(unsigned(IR(11 downto 8)))   when RegA1SelCmd = RegA1SelCmd_Rn else
                to_integer(unsigned(IR(7 downto 4)))    when RegA1SelCmd = RegA1SelCmd_Rm else
                R15                                     when RegA1SelCmd = RegA1SelCmd_R15 else
                R0;

    RegAxInSel <= to_integer(unsigned(IR(11 downto 8))) when RegAxInSelCmd = RegAxInSelCmd_Rn else
                  to_integer(unsigned(IR(7 downto 4)))  when RegAxInSelCmd = RegAxInSelCmd_Rm else
                  R15                                   when RegAxInSelCmd = RegAxInSelCmd_R15 else
                  R0;

    -- Control Unit Registers
    process (CLK)
    begin

        if rising_edge(CLK) then

            if RST = '1' then
                -- Since databus is 32-bits, the IR is the high 16 bits when the
                -- program address when is at an address that is a multiple of 4.
                -- When it's not a multiple of 4 them the IR is the low 16 bits.
                IR <= DB(31 downto 16) when UpdateIR_EX = '1' and AB(1 downto 0) = "00" else
                      DB(15 downto 0) when UpdateIR_EX = '1' and AB(1 downto 0) = "10" else
                      IR;

                -- Update status register accordingly
                if UpdateSR_EX = '1' then
                    SR <= (31 downto 1 => '0') & Tbit  when SRSel = SRSel_Tbit else
                          DB                           when SRSel = SRSel_DB   else
                          RegB                         when SRSel = SRSel_Reg  else
                          TempReg2                     when SRSel = SRSel_Tmp2 else
                          (others => 'X');
                end if;

                -- Update temporary register 1
                TempReg <= TempRegMuxOut when UpdateTempReg = '1' else TempReg;

                -- Update temporary register 2
                TempReg2 <= TempReg2MuxOut when UpdateTempReg2 = '1' else TempReg2;

                -- Set state of FSM
                CurrentState <= NextState when ForceNormalStateNext = '0' else Normal;

            else
                -- Reset to idle instruction (rising edge after reset)
                -- IR <= OpBoot;
                IR <= OpNOP;
                CurrentState <= Normal;
            end if;

        end if;
    end process;
    
    process (all)
    begin

        -- Add default values to prevent inferred latches during synthesis
        ALUOpASel <= unused;
        ALUOpBSel <= unused;
        FCmd <= (others => '-');
        CinCmd <= (others => '-');
        SCmd <= (others => '-');
        ALUCmd <= (others => '-');
        TbitOp <= (others => '-');
        UpdateSR <= '0';
        PAU_SrcSel <= PAU_AddrPC;
        PAU_OffsetSel <= PAU_OffsetWord;
        PAU_UpdatePC <= '1';
        PAU_PRSel <= PRSel_None;
        PAU_IncDecBit <= unused;
        PAU_PrePostSel <= MemUnit_POST;
        PAU_IncDecSel <= '1';
        DAU_SrcSel <= unused;
        DAU_OffsetSel <= unused;
        DAU_IncDecSel <= '-';
        DAU_IncDecBit <= unused;
        DAU_PrePostSel <= '-';
        DAU_GBRSel <= GBRSel_None;
        DAU_VBRSel <= VBRSel_None;
        RegInSelCmd <= RegInSelCmd_Rn;
        RegStore <= '0';
        RegASelCmd <= 0;
        RegBSelCmd <= 0;
        RegAxInSelCmd <= 0;
        RegAxStore <= '0';
        RegA1SelCmd <= 0;
        RegOpSel <= RegOpSel_None;
        RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
        RD <= '0';
        WR <= '1';
        ABOutSel <= ABOutSel_Prog;
        DBInMode <= 0;
        DBOutSel <= 0;
        DataAccessMode <= DataAccessMode_Word;
        NextState <= Normal;
        UpdateIR <= '1';
        UpdateTempReg <= '0';
        TempRegSel <= 0;
        TempReg2Sel <= 0;
        SRSel <= 0;
        UpdateTempReg2 <= '0';

    -- Instruction decoding (auto-generated)
    if std_match(IR, OpMOV_Imm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Signed;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_At_Disp_PC_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_At_Disp_PC_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOV_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_Rm_To_At_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_Rm_To_At_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_Rm_To_At_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_At_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_At_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_At_Rm_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_Rm_To_At_Dec_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 0;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_Rm_To_At_Dec_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 1;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_Rm_To_At_Dec_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_At_Rm_Inc_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rm;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_At_Rm_Inc_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 1;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rm;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_At_Rm_Inc_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rm;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_R0_To_At_Disp_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x1;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_R0_To_At_Disp_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_R0_To_At_Disp_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_At_Disp_Rm_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x1;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_At_Disp_Rm_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_At_Disp_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_Rm_To_At_R0_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_Rm_To_At_R0_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_Rm_To_At_R0_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_At_R0_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_At_R0_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_At_R0_Rm_To_Rn) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_R0_To_At_Disp_GBR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x1;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_R0_To_At_Disp_GBR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_R0_To_At_Disp_GBR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVB_At_Disp_GBR_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x1;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVW_At_Disp_GBR_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVL_At_Disp_GBR_To_R0) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Signed;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVA) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_R0;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rm;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_DataAddr;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpMOVT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Tbit;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSwapB) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SWAPB;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSwapW) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SWAPW;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpXTRCT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_XTRCT;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= DBInMode_Signed;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpADD_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_ADDER;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpADD_Imm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Signed;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_ADDER;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpADDC) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_CIN;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpADDV) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Overflow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_EQ_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Signed;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_EQ_RmRn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_HS) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_GE) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GEQ;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_HI) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_HI;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_GT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GT;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_PL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_Zero;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_PL;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_PZ) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_Zero;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_PZ;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCMP_STR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_STR;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpDT) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_ONE;
			CinCmd <= CinCmd_Zero;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpEXTS_B) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_EXTSB;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpEXTS_W) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_EXTSW;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpEXTU_B) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_EXTUB;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpEXTU_W) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_EXTUW;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpNEG) then
			ALUOpASel <= ALUOpASel_Zero;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpNEGC) then
			ALUOpASel <= ALUOpASel_Zero;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_CINBAR;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Borrow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSUB) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSUBC) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_CINBAR;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Borrow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSUBV) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Overflow;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpAND_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_AND;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpAND_Imm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpAND_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WriteBack;
			UpdateIR <= '0';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Result;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '1';
			TempReg2Sel <= TempReg2Sel_Result;
		elsif std_match(IR, OpNOT) then
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_NOTB;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpOR_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_OR;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpOR_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_OR;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpOR_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_OR;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WriteBack;
			UpdateIR <= '0';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Result;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '1';
			TempReg2Sel <= TempReg2Sel_Result;
		elsif std_match(IR, OpTAS_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_TASMask;
			FCmd <= FCmd_OR;
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_TAS;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WriteBack;
			UpdateIR <= '0';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Result;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '1';
			TempReg2Sel <= TempReg2Sel_Result;
		elsif std_match(IR, OpTST_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_AND;
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpTST_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpTST_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_AND;
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Result;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '1';
			TempReg2Sel <= TempReg2Sel_Result;
		elsif std_match(IR, OpXOR_Rm_Rn) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_XOR;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpXOR_Imm) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_XOR;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_R0;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpXOR_Imm_B) then
			ALUOpASel <= ALUOpASel_DB;
			ALUOpBSel <= ALUOpBSel_Imm_Unsigned;
			FCmd <= FCmd_XOR;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_R0;
			RegBSelCmd <= RegBSelCmd_R0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_R0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Unsigned;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WriteBack;
			UpdateIR <= '0';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Result;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '1';
			TempReg2Sel <= TempReg2Sel_Result;
		elsif std_match(IR, OpROTL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_ROL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpROTR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_ROR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpROTCL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_RLC;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpROTCR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_RRC;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHAL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_LSL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHAR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_ASR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLL) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_LSL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLR) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			SCmd <= SCmd_LSR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLL2) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SHLL2;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLR2) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SHLR2;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLL8) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SHLL8;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLR8) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SHLR8;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLL16) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SHLL16;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSHLR16) then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			FCmd <= FCmd_B;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '1';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_SHLR16;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBF) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when SR(0) = '0' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBFS) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot when SR(0)='0' else Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset8;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBT) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when SR(0) = '1' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBTS) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot when SR(0)='1' else Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset8;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBRA) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset12;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBRAF) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBSR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_PC;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_Offset12;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBSRF) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_PC;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlot;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpJMP) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlotDirect;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpJSR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_PC;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxStore <= '0';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlotDirect;
			UpdateIR <= '1';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpRTS) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= BranchSlotRet;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= TempRegSel_RegB;
			SRSel <= SRSel_Tbit;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpCLRT) then
			FCmd <= FCmd_ONE;
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDC_Rm_To_SR) then
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= SRSel_Reg;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDC_Rm_To_GBR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_GBRSel <= GBRSel_Reg;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDC_Rm_To_VBR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_Reg;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_SR) then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= SRSel_DB;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_GBR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_DB;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_VBR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_DB;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDS_Rm_To_PR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_Reg;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= RegASelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpLDSL_At_Rm_Inc_To_PR) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_DB;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rm;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSLEEP) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Sleep;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpNOP) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpRTE) then
			UpdateSR <= '0';
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= RegASelCmd_Rn;
			RegBSelCmd <= RegBSelCmd_Rn;
			RegAxInSelCmd <= RegAxInSelCmd_R15;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_R15;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= RTE_PopSR;
			UpdateIR <= '0';
			UpdateTempReg <= '1';
			TempRegSel <= TempRegSel_DataBus;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSETT) then
			FCmd <= FCmd_ZERO;
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTC_SR_To_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_SR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTC_GBR_To_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_GBR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTC_VBR_To_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_VBR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTCL_SR_To_At_Dec_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_SR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTCL_GBR_To_At_Dec_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_GBR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTCL_VBR_To_At_Dec_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_VBR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTS_PR_To_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_PR;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpSTSL_PR_To_At_Dec_Rn) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_Rn;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_Rn;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_PR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpTRAPA) then
			UpdateSR <= '0';
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= RegAxInSelCmd_R15;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_R15;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= DBOutSel_SR;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= TRAPA_PushPC;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		elsif std_match(IR, OpBoot) then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrDB;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			PAU_PrePostSel <= MemUnit_POST;
			PAU_IncDecSel <= '1';
			DAU_SrcSel <= DAU_AddrZero;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegInSelCmd <= RegInSelCmd_Rn;
			RegStore <= '0';
			RegASelCmd <= 0;
			RegBSelCmd <= 0;
			RegAxInSelCmd <= 0;
			RegAxStore <= '0';
			RegA1SelCmd <= 0;
			RegOpSel <= RegOpSel_None;
			RegAxInDataSel <= 0;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= 0;
			DBOutSel <= 0;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= BootReadSP;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			TempRegSel <= 0;
			SRSel <= 0;
			UpdateTempReg2 <= '0';
		end if;

		-- State Decoding Autogen
		if CurrentState = WaitForFetch then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			DAU_GBRSel <= 0;
			DAU_VBRSel <= 0;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = Sleep then
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			DAU_GBRSel <= 0;
			DAU_VBRSel <= 0;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RD <= '1';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Sleep;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = BranchSlot then
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_TempReg;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 1;
			PAU_PrePostSel <= MemUnit_PRE;
			PAU_IncDecSel <= MemUnit_DEC;
		elsif CurrentState = BranchSlotRet then
			PAU_SrcSel <= PAU_AddrPR;
			PAU_OffsetSel <= PAU_OffsetLong;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = BranchSlotDirect then
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_TempReg;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = BootReadSP then
			ALUOpASel <= ALUOpASel_DB;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_UpdatePC <= '0';
			PAU_PRSel <= PRSel_None;
			DAU_SrcSel <= DAU_AddrZero;
			DAU_OffsetSel <= DAU_OffsetLong;
			DAU_PrePostSel <= MemUnit_POST;
			RegInSelCmd <= RegInSelCmd_R15;
			RegStore <= '1';
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= BootWaitForFetch;
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_PRE;
		elsif CurrentState = BootWaitForFetch then
			ALUOpASel <= ALUOpASel_RegA;
			ALUOpBSel <= ALUOpBSel_RegB;
			UpdateSR <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			DAU_GBRSel <= 0;
			DAU_VBRSel <= 0;
			RegStore <= '0';
			RegAxStore <= '0';
			RegOpSel <= RegOpSel_None;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = WriteBack then
			ALUOpASel <= ALUOpASel_TempReg;
			FCmd <= FCmd_A;
			ALUCmd <= ALUCmd_FBLOCK;
			UpdateSR <= '0';
			PAU_UpdatePC <= '0';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegStore <= '0';
			RegAxStore <= '0';
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBOutSel <= DBOutSel_Result;
			DataAccessMode <= DataAccessMode_Byte;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 0;
			PAU_PrePostSel <= MemUnit_POST;
		elsif CurrentState = TRAPA_PushPC then
			PAU_UpdatePC <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegStore <= '0';
			RegAxInSelCmd <= RegAxInSelCmd_R15;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_R15;
			RD <= '1';
			WR <= '0';
			ABOutSel <= ABOutSel_Data;
			DBOutSel <= DBOutSel_PC;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= TRAPA_ReadVector;
			UpdateIR <= '0';
		elsif CurrentState = TRAPA_ReadVector then
			PAU_SrcSel <= PAU_AddrDB;
			PAU_OffsetSel <= PAU_OffsetZero;
			PAU_UpdatePC <= '1';
			DAU_SrcSel <= DAU_AddrVBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegStore <= '0';
			RegAxInSelCmd <= RegAxInSelCmd_R15;
			RegAxStore <= '0';
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DBInMode <= DBInMode_Unsigned;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= WaitForFetch;
			UpdateIR <= '0';
		elsif CurrentState = RTE_PopSR then
			PAU_UpdatePC <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_GBRSel <= GBRSel_None;
			DAU_VBRSel <= VBRSel_None;
			RegStore <= '0';
			RegAxInSelCmd <= RegAxInSelCmd_R15;
			RegAxInDataSel <= RegAxInDataSel_AddrIDOut;
			RegAxStore <= '1';
			RegA1SelCmd <= RegA1SelCmd_R15;
			RD <= '0';
			WR <= '1';
			ABOutSel <= ABOutSel_Data;
			DataAccessMode <= DataAccessMode_Long;
			NextState <= RTE_Slot;
			UpdateIR <= '0';
			UpdateTempReg <= '0';
			UpdateTempReg2 <= '1';
			TempReg2Sel <= TempReg2Sel_DB;
			SRSel <= SRSel_Tmp2;
		elsif CurrentState = RTE_Slot then
			UpdateSR <= '1';
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_TempReg;
			PAU_UpdatePC <= '1';
			PAU_PRSel <= PRSel_None;
			RegStore <= '0';
			RegAxInSelCmd <= RegAxInSelCmd_R15;
			RegAxStore <= '0';
			ABOutSel <= ABOutSel_Prog;
			DataAccessMode <= DataAccessMode_Word;
			NextState <= Normal;
			UpdateIR <= '1';
			UpdateTempReg <= '0';
			PAU_IncDecBit <= 1;
			PAU_PrePostSel <= MemUnit_PRE;
			PAU_IncDecSel <= MemUnit_INC;
			SRSel <= SRSel_Tmp2;
		end if;


    -- end of auto-generated code (continue process)
        
    end process;


end behavioral;
