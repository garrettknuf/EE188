----------------------------------------------------------------------------
--
--  SH-2 Control Unit
--
--  This is an implementation of 
--
--  Entities included are:
--    
--
--  Revision History:
--     18 April 2025    Garrett Knuf    Initial revision.
--
----------------------------------------------------------------------------

--
-- Package containing constants for the control unit.
--

library ieee;
use ieee.std_logic_1164.all;
use work.GenericConstants.all;

package CUConstants is

    -- Data Transfer Instructions (Table 5.3)
    constant OpMOV_Imm_To_Rn          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "1110------------";
    constant OpMOVW_Disp_PC_To_Rn     : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "1001------------";
    constant OpMOVL_Disp_PC_To_Rn     : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "1101------------";
    constant OpMOV_Rm_To_Rn           : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0011";
    constant OpMOVB_Rm_To_At_Rn       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------0000";
    constant OpMOVW_Rm_To_At_Rn       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------0001";
    constant OpMOVL_Rm_To_At_Rn       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------0010";
    constant OpMOVB_At_Rm_To_Rn       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0000";
    constant OpMOVW_At_Rm_To_Rn       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0001";
    constant OpMOVL_At_Rm_Rn          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0010";
    constant OpMOVB_Rm_To_At_Dec_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------0000";
    constant OpMOVW_Rm_To_At_Dec_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------0001";
    constant OpMOVL_Rm_To_At_Dec_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------0010";
    constant OpMOVB_At_Rm_Inc_To_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0100";
    constant OpMOVW_At_Rm_Inc_To_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0101";
    constant OpMOVL_At_Rm_Inc_To_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0110";
    constant OpMOVB_R0_To_At_Disp_Rn  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10000000--------";
    constant OpMOVW_R0_To_At_Disp_Rn  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10000001--------";
    constant OpMOVL_R0_To_At_Disp_Rn  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0001------------";
    constant OpMOVB_At_Disp_Rm_To_R0  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10000100--------";
    constant OpMOVW_At_Disp_Rm_To_R0  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10000101--------";
    constant OpMOVL_At_Disp_Rm_To_Rn  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0101------------";
    constant OpMOVB_Rm_To_At_R0_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000--------0100";
    constant OpMOVW_Rm_To_At_R0_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000--------0101";
    constant OpMOVL_Rm_To_At_R0_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000--------0100";
    constant OpMOVB_At_R0_Rm_To_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000--------1100";
    constant OpMOVW_At_R0_Rm_To_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000--------1101";
    constant OpMOVL_At_R0_Rm_To_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000--------1110";
    constant OpMOVB_R0_To_At_Disp_GBR : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000000--------";
    constant OpMOVW_R0_To_At_Disp_GBR : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000001--------";
    constant OpMOVL_R0_To_At_Disp_GBR : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000010--------";
    constant OpMOVB_At_Disp_GBR_To_R0 : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000100--------";
    constant OpMOVW_At_Disp_GBR_To_R0 : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000101--------";
    constant OpMOVL_At_Disp_GBR_To_R0 : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000110--------";
    constant OpMOVA                   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000111--------";
    constant OpMOVT                   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00101001";
    constant OpSwapB                  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1000";
    constant OpSwapW                  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1001";
    constant OpXTRCT                  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------1101";

    -- Arithmetic Instructions (Table 5.4)
    constant OpADD_Rm_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------1100";
    constant OpADD_Imm_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0111------------";
    constant OpADDC         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------1110";
    constant OpADDV         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------1111";
    constant OpCMP_EQ_Imm   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10001000--------";
    constant OpCMP_EQ_RmRn  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------0000";
    constant OpCMP_HS       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------0010";
    constant OpCMP_GE       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------0011";
    constant OpCMP_HI       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------0110";
    constant OpCMP_GT       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------0111";
    constant OpCMP_PL       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00010101";
    constant OpCMP_PZ       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00010001";
    constant OpCMP_STR      : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------1100";
    -- TODO: DIV1
    -- TODO: DIV0S
    -- TODO: DIV0U
    -- TODO: DMULS.L
    -- TODO: DMULU.L
    constant OpCMP_DT       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00010000";
    constant OpEXTS_B       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1110";
    constant OpEXTS_W       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1111";
    constant OpEXTU_B       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1100";
    constant OpEXTU_W       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1101";
    -- TODO: MAC.L
    -- TODO: MAC.W
    -- TODO: MUL.L
    -- TODO: MULS.W
    -- TODO: MULU.W
    constant OpNEG          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1011";
    constant OpNEGC         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------1010";
    constant OpSUB          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------1000";
    constant OpSUBC         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------1010";
    constant OpSUBV         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0011--------1011";

    -- Logic Operation Instructions (Table 5.5)
    constant OpAND_Rm_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------1001";
    constant OpAND_Imm_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001001--------";
    constant OpAND_Imm_B    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001101--------";
    constant OpNOT          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0110--------0111";
    constant OpOR_Rm_Rn     : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------1011";
    constant OpOR_Imm       : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001011--------";
    constant OpOR_Imm_B     : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001011--------";
    constant OpTAS_B        : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00011011";
    constant OpTST_Rm_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------1000";
    constant OpTST_Imm      : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001000--------";
    constant OpTST_Imm_B    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001100--------";
    constant OpXOR_Rm_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0010--------1010";
    constant OpXOR_Imm      : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001010--------";
    constant OpXOR_Imm_B    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11001110--------";

    -- Shift Instructions (Table 5.6)
    constant OpROTL         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00000100";
    constant OpROTR         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00000101";
    constant OpROTCL        : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100100";
    constant OpROTCR        : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100101";
    constant OpSHAL         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100000";
    constant OpSHAR         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100001";
    constant OpSHLL         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00000000";
    constant OpSHLR         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00000001";
    -- TODO: SHLL2
    -- TODO: SHLR2
    -- TODO: SHLL8
    -- TODO: SHLR8
    -- TODO: SHLL16
    -- TODO: SHLR16

    -- Branch Instructions (Table 5.7)
    constant OpBF           : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10001011--------";
    constant OpBFS          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10001111--------";
    constant OpBT           : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10001001--------";
    constant OpBTS          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "10001101--------";
    constant OpBRA          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "1010------------";
    constant OpBRAF         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00100011";
    constant OpBSR          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "1011------------";
    constant OpBSRF         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00000011";
    constant OpJMP          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00101011";
    constant OpJSR          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00001011";
    constant OpRTS          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000000000001011";

    -- System Control Instructions (Table 5.8)
    constant OpCLRT                  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000000000001000";
    -- TODO: CLRMAC
    constant OpLDC_Rm_To_SR          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00001110";
    constant OpLDC_Rm_To_GBR         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00011110";
    constant OpLDC_Rm_To_VBR         : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00101110";
    constant OpLDCL_At_Rm_Inc_To_SR  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00000111";
    constant OpLDCL_At_Rm_Inc_To_GBR : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00010111";
    constant OpLDCL_At_Rm_Inc_To_VBR : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100111";
    -- TODO: LDS Rm, MACH
    -- TODO: LDS Rm, MACL
    constant OpLDS_Rm_To_PR          : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00101010";
    -- TODO: LDS.L @Rm+, MACH
    -- TODO: LDS.L @Rm+, MACL
    constant OpLDSL_At_Rm_Inc_To_PR  : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00101010";
    constant NOP                     : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000000000001001";
    constant RTE                     : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000000000101011";
    -- TODO: Sleep
    constant STC_SR_To_Rn            : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00000010";
    constant STC_GBR_To_Rn           : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00010010";
    constant STC_VBR_To_Rn           : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00100010";
    constant STCL_SR_To_At_Dec_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00000011";
    constant STCL_GBR_To_At_Dec_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00010011";
    constant STCL_VBR_To_At_Dec_Rn   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100011";
    -- TODO: STS MACH, Rn
    -- TODO: STS MACL, Rn
    -- TODO: STS MACH, Rn
    constant STS_PR_To_Rn            : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0000----00101010";
    -- TODO: STSL MACH, @-Rn
    -- TODO: STSL MACL, @-Rn
    constant STSL_PR_To_At_Dec_Rn    : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "0100----00100010";
    constant TRAPA                   : std_logic_vector(DATA_BUS_SIZE-1 downto 0) := "11000011--------";


    constant ALUOpACmd_RegA  : std_logic_vector(1 downto 0) := "00";

    constant ALUOPBCMD_SrcCnt : integer := 2;
    constant ALUOpBCmd_RegB   : integer range ALUOPBCMD_SrcCnt - 1 downto 0 := 0;
    constant ALUOpBCmd_IR_Imm : integer range ALUOPBCMD_SrcCnt - 1 downto 0 := 1;

    constant BusCmd_Prog := std_logic := '0';
    constant BusCmd_Data := std_logic := '1';
    



end package;


--
--
--
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.GenericConstants.all;
use work.CUConstants.all;
use work.ALUConstants.all;
use work.TbitConstants.all;
use work.DAUConstants.all;
use work.PAUConstants.all;
use work.RegArrayConstants.all;
use work.StatusRegConstants.all;

entity CU is

    port (
        -- CU Input Signals
        CLK     : in    std_logic;
        DB      : in    std_logic_vector(DATA_BUS_SIZE - 1 downto 0);
        SR      : in    std_logic_vector(REG_SIZE - 1 downto 0);

        -- ALU Control Signals
        ALUOpACmd   : out     std_logic_vector(1 downto 0);
        ALUOpBCmd   : out     std_logic_vector(1 downto 0);                          
        FCmd        : out     std_logic_vector(3 downto 0);            
        CinCmd      : out     std_logic_vector(1 downto 0);            
        SCmd        : out     std_logic_vector(2 downto 0);            
        ALUCmd      : out     std_logic_vector(1 downto 0);
        TbitOp      : out     integer range Tbit_Src_Cnt - 1 downto 0; 

        -- StatusReg Control Signals
        UpdateTbit  : out   std_logic

        -- RegArray Control Signals
        RegInSel   : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegStore   : out   std_logic;
        RegASel    : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegBSel    : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegAxInSel : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegAxStore : out   std_logic;
        RegA1Sel   : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegA2Sel   : out   integer  range REGARRAY_RegCnt - 1 downto 0;
        RegOpSel   : out   integer  range REGOp_SrcCnt - 1 downto 0;
        
        -- DAU Control Signals
        DAU_SrcSel      : out   integer range DAU_SRC_CNT - 1 downto 0;
        DAU_OffsetSel   : out   integer range DAU_OFFSET_CNT - 1 downto 0;
        DAU_IncDecSel   : out   std_logic;
        DAU_IncDecBit   : out   integer range 2 downto 0;
        DAU_PrePostSel  : out   std_logic;
        DAU_LoadGBR     : out   std_logic;

        -- PAU Control Signals
        PAU_SrcSel      : out   integer range PAU_SRC_CNT - 1 downto 0;
        PAU_OffsetSel   : out   integer range PAU_OFFSET_CNT - 1 downto 0;
        PAU_UpdatePC    : out   std_logic;
        PAU_UpdatePR    : out   std_logic;

    );

end CU;

architecture behavioral of CU is

    signal IR : std_logic_vector(DATA_BUS_SIZE-1 downto 0);

begin

    -- Control Unit FSM
    process (CLK)
    begin

        if rising_edge(CLK) then

            -- Temporary only reading from memory (fetch)
            IR <= DB;

        end if;

    end process;

    -- Instruction decoding (auto-generated)
    process (all)
	begin
		if std_match(IR, OpMOV_Imm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpMOVW_Disp_PC_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVL_Disp_PC_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOV_Rm_To_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpMOVB_Rm_To_At_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVW_Rm_To_At_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVL_Rm_To_At_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVB_At_Rm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVW_At_Rm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVL_At_Rm_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVB_Rm_To_At_Dec_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVW_Rm_To_At_Dec_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= '1';
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVL_Rm_To_At_Dec_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVB_At_Rm_Inc_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVW_At_Rm_Inc_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= '1';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVL_At_Rm_Inc_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVB_R0_To_At_Disp_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_R0;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVW_R0_To_At_Disp_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_R0;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVL_R0_To_At_Disp_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x3;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_R0;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVB_At_Disp_Rm_To_R0) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= R0;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVW_At_Disp_Rm_To_R0) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= R0;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVL_At_Disp_Rm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_Offset4x3;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVB_Rm_To_At_R0_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVW_Rm_To_At_R0_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVL_Rm_To_At_R0_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rn;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVB_At_R0_Rm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVW_At_R0_Rm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVL_At_R0_Rm_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetR0;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVB_R0_To_At_Disp_GBR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_R0;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rm;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVW_R0_To_At_Disp_GBR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_R0;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rm;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVL_R0_To_At_Disp_GBR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_R0;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rm;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, OpMOVB_At_Disp_GBR_To_R0) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x1;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= R0;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVW_At_Disp_GBR_To_R0) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x2;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= R0;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVL_At_Disp_GBR_To_R0) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrGBR;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= R0;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVA) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrPC;
			DAU_OffsetSel <= DAU_Offset8x4;
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= R0;
			RegStore <= '1';
			RegASel <= RegASel_Rm;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rm;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpMOVT) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= RegAxInSel_Rm;
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSwapB) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSwapW) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpXTRCT) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpADD_Rm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpADD_Imm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpADDC) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Carry;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpADDV) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_B;
			CinCmd <= CinCmd_Zero;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Overflow;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_EQ_Imm) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_EQ_RmRn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_HS) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GEQ;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_GE) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GEQ;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_HI) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_HI;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_GT) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_GT;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_PL) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_Zero;
			CinCmd <= CinCmd_Zero;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_PL;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_PZ) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_Zero;
			CinCmd <= CinCmd_Zero;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_PZ;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_STR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_STR;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCMP_DT) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_Zero;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpEXTS_B) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpEXTS_W) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpEXTU_B) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpEXTU_W) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_A;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpNEG) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_NOTA;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpNEGC) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_NOTA;
			CinCmd <= CinCmd_Borrow;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Borrow;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSUB) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSUBC) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_Borrow;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Borrow;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSUBV) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOTB;
			CinCmd <= CinCmd_One;
			SCmd <= '-';
			ALUCmd <= ALUCmd_ADDER;
			TbitOp <= Tbit_Overflow;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpAND_Rm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_AND;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpAND_Imm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_AND;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpAND_Imm_B) then
			ALUOpACmd <= ALUOpACmd_DB;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_AND;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForRead;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpNOT) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_NOT;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpOR_Rm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_OR;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpOR_Imm) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_OR;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpOR_Imm_B) then
			ALUOpACmd <= ALUOpACmd_DB;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_OR;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForRead;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpTAS_B) then
			ALUOpACmd <= ALUOpACmd_DB;
			ALUOpBCmd <= '-';
			FCmd <= FCmd_ONES;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForRead;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpTST_Rm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_AND;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpTST_Imm) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_AND;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '0';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpTST_Imm_B) then
			ALUOpACmd <= ALUOpACmd_DB;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_AND;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForRead;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpXOR_Rm_Rn) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_RegB;
			FCmd <= FCmd_XOR;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= RegBSel_Rm;
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpXOR_Imm) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_XOR;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpXOR_Imm_B) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= ALUOpBCmd_Imm;
			FCmd <= FCmd_XOR;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForRead;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpROTL) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_ROL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpROTR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_ROR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpROTCL) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_RLC;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpROTCR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_RRC;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHAL) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHAR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_ASR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLL) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSL;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLR) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSR;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= Tbit_Carry;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLL2) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSL2;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLR2) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSR2;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLL8) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSL8;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLR8) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSR8;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLL16) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSL16;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpSHLR16) then
			ALUOpACmd <= ALUOpACmd_RegA;
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= SCmd_LSR16;
			ALUCmd <= ALUCmd_SHIFT;
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= RegInSel_Rn;
			RegStore <= '1';
			RegASel <= RegASel_Rn;
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBF) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when Tbit = '0' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= BranchSlot when Tbit = '0' else Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBFS) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when Tbit = '0' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= BranchSlot when Tbit = '0' else Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBT) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when Tbit = '1' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= BranchSlot when Tbit = '1' else Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBTS) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset8 when Tbit = '1' else PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= BranchSlot when Tbit = '1' else Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBRA) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset12;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBRAF) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetReg;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= RegA1Sel_IR_11_8;
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBSR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_Offset12;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '1';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpBSRF) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetReg;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '1';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= RegA1Sel_IR_11_8;
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpJMP) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_OffsetReg;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= RegA1Sel_IR_11_8;
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpJSR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_OffsetReg;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '1';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= RegA1Sel_IR_11_8;
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpRTS) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrZero;
			PAU_OffsetSel <= PAU_OffsetPR;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '-';
			RegStore <= '0';
			RegASel <= '-';
			RegBSel <= '-';
			RegAxInSel <= '-';
			RegAxStore <= '0';
			RegA1Sel <= '-';
			RegA2Sel <= '-';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpCLRT) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= FCmd_ONE;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpLDC_Rm_To_SR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpLDC_Rm_To_GBR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '1';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpLDC_Rm_To_VBR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_SR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '1';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForReadPostInc;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_GBR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '1';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForReadPostInc;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpLDCL_At_Rm_Inc_To_VBR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= WaitForReadPostInc;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, OpLDS_Rm_To_PR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= nan;
			PAU_OffsetSel <= nan;
			PAU_UpdatePC <= nan;
			PAU_UpdatePR <= nan;
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, OpLDSL_At_Rm_Inc_To_PR) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '1';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_INC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_POST;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '1';
			WR <= '0';
		elsif std_match(IR, NOP) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, RTE) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '1';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '1';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= RTE_Init;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, SETT) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= FCmd_ZERO;
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= ALUCmd_FBLOCK;
			TbitOp <= Tbit_Zero;
			UpdateTbit <= '1';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, STC_SR_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, STC_GBR_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, STC_VBR_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, STCL_SR_To_At_Dec_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, STCL_GBR_To_At_Dec_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, STCL_VBR_To_At_Dec_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Fetch;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, STS_PR_To_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '-';
			DAU_OffsetSel <= '-';
			DAU_IncDecSel <= '-';
			DAU_IncDecBit <= '-';
			DAU_PrePostSel <= '-';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '0';
		elsif std_match(IR, STSL_PR_To_At_Dec_Rn) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= PAU_AddrPC;
			PAU_OffsetSel <= PAU_OffsetWord;
			PAU_UpdatePC <= '1';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= DAU_AddrRn;
			DAU_OffsetSel <= DAU_OffsetZero;
			DAU_IncDecSel <= MemUnit_DEC;
			DAU_IncDecBit <= 2;
			DAU_PrePostSel <= MemUnit_PRE;
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= Idle;
			RD <= '0';
			WR <= '1';
		elsif std_match(IR, TRAPA) then
			ALUOpACmd <= '-';
			ALUOpBCmd <= '-';
			FCmd <= '-';
			CinCmd <= '-';
			SCmd <= '-';
			ALUCmd <= '-';
			TbitOp <= '-';
			UpdateTbit <= '0';
			PAU_SrcSel <= '-';
			PAU_OffsetSel <= '-';
			PAU_UpdatePC <= '0';
			PAU_UpdatePR <= '0';
			DAU_SrcSel <= '0';
			DAU_OffsetSel <= '0';
			DAU_IncDecSel <= '0';
			DAU_IncDecBit <= '0';
			DAU_PrePostSel <= '0';
			DAU_LoadGBR <= '0';
			RegInSel <= '0';
			RegStore <= '0';
			RegASel <= '0';
			RegBSel <= '0';
			RegAxInSel <= '0';
			RegAxStore <= '0';
			RegA1Sel <= '0';
			RegA2Sel <= '0';
			RegOpSel <= '0';
			NextState <= TRAPA_Init;
			RD <= '1';
			WR <= '0';
		end if;
	 end process;


end behavioral;
